//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-3
//Part Number: GW2AR-LV18EQ144C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Thu May 09 15:00:13 2024

module table_FONT (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [16:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [0:0] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [0:0] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [0:0] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [0:0] prom_inst_7_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_0.INIT = 16'h0002;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_1.INIT = 16'h0008;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_2.INIT = 16'h0020;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_3.INIT = 16'h0080;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_4.INIT = 16'h0200;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_5.INIT = 16'h0800;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_6.INIT = 16'h2000;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_7.INIT = 16'h8000;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0001800000018000078001E0078001E000000000000000000000FFFFFFFF0000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000C30000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h0180018001800000018001800180000000000180000000000000000000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h0003C0000003C0001F8001F81F8001F800000000000000000000FFFF80010000;
defparam prom_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'h1000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h0000000000000008000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h00000000000000000000000006E0000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0180018001800000018001800180000000000180000000000000000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h1803C0181803C0183000001C3000001C003F0000003F00000000FFFF80010000;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h1000000000000000000000000000000000000000000001000440000000000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0000000000000008000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000040;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h00000000000000000000000003C0000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h0180018001800000018001800180000000000180000000000000000000000000;
defparam prom_inst_0.INIT_RAM_30 = 256'h3C03C03C3C03C03C600000066000000600E1C00000E1C0000040FFFF80010000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h1000000000000000000000000000000000000000004001000440000001800000;
defparam prom_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000380038000001C000000000003C003C001000380;
defparam prom_inst_0.INIT_RAM_34 = 256'h00000000000000000000000000000000000000000000000000000000000003C0;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000008000000018000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h00000000000000000000000000000000000000000000000000000000000000C0;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0180018001800000018001800180000000000180000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h3E03C07C3E03C07C4001800640018006018060000180600001B0FFFF80010000;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h08000000000003C0000001800010080003C0000001B001000440071C01800000;
defparam prom_inst_1.INIT_RAM_03 = 256'h00000000000000000000000007C007E01FF83F000FF0060007E007E001C007E0;
defparam prom_inst_1.INIT_RAM_04 = 256'h00000000000000000000000000000000000000000000000000000000000007E0;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000018001F000100F0000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000001C00007F0000001E000000000E00000080;
defparam prom_inst_1.INIT_RAM_07 = 256'h0000000000E00100060000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0A = 256'h0000000000000000000000000810000000000000000000000000000010000000;
defparam prom_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000001E00000000000000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C00080000000;
defparam prom_inst_1.INIT_RAM_0F = 256'h018001800180000001800180018000000000018000000000000000000000FFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'h1F03C0F81F03C0F8C0018003C001800303003000030030000110FFFF80010000;
defparam prom_inst_1.INIT_RAM_11 = 256'h3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C;
defparam prom_inst_1.INIT_RAM_12 = 256'h080000000000038000000180003008000380000001100FC00440063801803C7C;
defparam prom_inst_1.INIT_RAM_13 = 256'h07E0000000000000000000000C600C3010080180001005000C300C3001F00C20;
defparam prom_inst_1.INIT_RAM_14 = 256'h03C07C0EF00E01FC7C7EFFC01FF83C7C27C07FFC3FFE03FC27C003FE00FC0C20;
defparam prom_inst_1.INIT_RAM_15 = 256'h000001800100001001001FF8783E783E7C3EF83F7C3E3FFC17C003FE03C007F8;
defparam prom_inst_1.INIT_RAM_16 = 256'h00000000000000F8000000000000001C00006180000018000000000800000180;
defparam prom_inst_1.INIT_RAM_17 = 256'h3C7C000000800100030000000000000000000000000000200000000000000000;
defparam prom_inst_1.INIT_RAM_18 = 256'h7FFE03C03C7CF00E7FF8707C703E703E07C443C23FFE7FF87FFC03FE3FFE01F8;
defparam prom_inst_1.INIT_RAM_19 = 256'h7FC01E1F07E4007EF81F00FF73DF73DF7C3E7C3E783E03C0F81E3FFC27C007F8;
defparam prom_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000810000000000000000000000000000018000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000001E00000000000000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h0003C0003C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'h018001800180000001800180018000000000018000003C7C3C7C3C7C0000FFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'h0F8181F00F8181F0C0018003C001800306001800060018000208FFFF80010000;
defparam prom_inst_1.INIT_RAM_21 = 256'h3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C;
defparam prom_inst_1.INIT_RAM_22 = 256'h08000000000003800000018000200C000380000002081E6004400E3001803C7C;
defparam prom_inst_1.INIT_RAM_23 = 256'h0E700000000000000000000008300810100800C0001005000818081801180830;
defparam prom_inst_1.INIT_RAM_24 = 256'h0E607C1EF00E03FC7C7EFFC01FF83C7C3C607FFC3FFE0FFC2E600FFE00FC0810;
defparam prom_inst_1.INIT_RAM_25 = 256'h000002C00100003001001FF87C3E7C3EFC3FFC3F7C7E3FFC1E700FFE0E601FFC;
defparam prom_inst_1.INIT_RAM_26 = 256'h00000000000000F8000000000000001800000080000018000000000800000300;
defparam prom_inst_1.INIT_RAM_27 = 256'h3C7C000001800100010000000000000000000000000000200000000000000000;
defparam prom_inst_1.INIT_RAM_28 = 256'h7FFE0E603C7CF00E7FF8787CF07EF07E0C64E3C63FFE7FF87FFC0FFE3FFE01F8;
defparam prom_inst_1.INIT_RAM_29 = 256'h7FE0331F0E74007EF83F01FFFBDFFBDF7E3E7E7E7C3E07E0F83E3FFC2E601FFC;
defparam prom_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000C3000000000000000000000000000000FE00000;
defparam prom_inst_1.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000001000000000000000000;
defparam prom_inst_1.INIT_RAM_2C = 256'h0003C0003C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_1.INIT_RAM_2F = 256'h018001800180000001800180018000000000018000003C7C3C7C3C7C0000FFFF;
defparam prom_inst_1.INIT_RAM_30 = 256'h07C7E3E007C7E3E0C0018003C0018003060C1800060018000208FFFF80010000;
defparam prom_inst_1.INIT_RAM_31 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_1.INIT_RAM_32 = 256'h04000000000001800100018000200400018007800208183004400C3001801018;
defparam prom_inst_1.INIT_RAM_33 = 256'h0810000C00003000000000001810181018080040001005801000180801000810;
defparam prom_inst_1.INIT_RAM_34 = 256'h1810301830140020101808000100101830304010301818103810180801C00810;
defparam prom_inst_1.INIT_RAM_35 = 256'h0000024001000020010010081008100820042004100821041810081818101020;
defparam prom_inst_1.INIT_RAM_36 = 256'h00000000000000700000000001800018000000C0000018000000000800000200;
defparam prom_inst_1.INIT_RAM_37 = 256'h1018000001000100010000000000000000000000000000200000000000000000;
defparam prom_inst_1.INIT_RAM_38 = 256'h10081810101830141020481018081808181CB10A301810204020180830080380;
defparam prom_inst_1.INIT_RAM_39 = 256'h10306184181C000820040021210421041008100810080100200C210438101020;
defparam prom_inst_1.INIT_RAM_3A = 256'h00000000000000000000000006E0000000000000000000000000000007F00000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000001000000000000000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_1.INIT_RAM_3D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_1.INIT_RAM_3F = 256'h018001800180000001800180018000000000018000001018101810180000FFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h03DFFBC003DFFBC0C007E003C007E0030C0C0C000C000C000208FFFF80010000;
defparam prom_inst_2.INIT_RAM_01 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_2.INIT_RAM_02 = 256'h04000000000001800100118800600400018007C00208181004400C7001801018;
defparam prom_inst_2.INIT_RAM_03 = 256'h1810001800001800000000001010101808000020001004801000100801001810;
defparam prom_inst_2.INIT_RAM_04 = 256'h1018303838140020081808000100101820184010301810103018100801200818;
defparam prom_inst_2.INIT_RAM_05 = 256'h0000046001000020010008081818181820042004100821041018181810182020;
defparam prom_inst_2.INIT_RAM_06 = 256'h00000000000000600000000003C0001800000040000018000000000800000000;
defparam prom_inst_2.INIT_RAM_07 = 256'h1018000001000100010000000000000000000000000000200000000000000000;
defparam prom_inst_2.INIT_RAM_08 = 256'h100810181018381410204C1018081808300C910A301810204020100830080240;
defparam prom_inst_2.INIT_RAM_09 = 256'h10184084100C0008200400212104210410081008181801003008210430182020;
defparam prom_inst_2.INIT_RAM_0A = 256'h00000000000000000000000003C0000000000000000000000000000000180000;
defparam prom_inst_2.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000001000000000000000000;
defparam prom_inst_2.INIT_RAM_0C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_2.INIT_RAM_0D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_2.INIT_RAM_0E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'h018001800180000001800180018000000000018000001018101810180000FFFF;
defparam prom_inst_2.INIT_RAM_10 = 256'h01FFFF8001FFFF80001C3800001C38000C0C0C000C000C000208FFFF80010000;
defparam prom_inst_2.INIT_RAM_11 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_2.INIT_RAM_12 = 256'h040000000000018001001DB80040060001800260020808100440186001801018;
defparam prom_inst_2.INIT_RAM_13 = 256'h1010003000000C00000000001010100808000020001004801000100801001018;
defparam prom_inst_2.INIT_RAM_14 = 256'h30083028281400200C1808000100101820084010301820102008100801200808;
defparam prom_inst_2.INIT_RAM_15 = 256'h00000C2001000060010008080810081020042008100821041008101830082020;
defparam prom_inst_2.INIT_RAM_16 = 256'h00000000000000600000000003C0001800000040000018000000000800000000;
defparam prom_inst_2.INIT_RAM_17 = 256'h1018000001000100010000000000000000000000000000200000000000000000;
defparam prom_inst_2.INIT_RAM_18 = 256'h1008300810182814102044101C081C08200C991A301810204020100830080240;
defparam prom_inst_2.INIT_RAM_19 = 256'h1008C0443004000820040021210421041008100808100FF01018210420082020;
defparam prom_inst_2.INIT_RAM_1A = 256'h00000000000000000000000000000000000000000000000000000000000C0000;
defparam prom_inst_2.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000001000000000000000000;
defparam prom_inst_2.INIT_RAM_1C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_2.INIT_RAM_1D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_2.INIT_RAM_1E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_2.INIT_RAM_1F = 256'h018001800180000001800180018000000000018000001018101810180000FFFF;
defparam prom_inst_2.INIT_RAM_20 = 256'h007FFE00007E7E0000300C0000300C00080C0400080004000108FFFF80010000;
defparam prom_inst_2.INIT_RAM_21 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_2.INIT_RAM_22 = 256'h0200000000000180010007E00040060001800020010800100440186001801018;
defparam prom_inst_2.INIT_RAM_23 = 256'h100000E000000600000000001010101808000010001004401000100001001008;
defparam prom_inst_2.INIT_RAM_24 = 256'h200C3028283400200618080001001018200C401030182010200C300801200808;
defparam prom_inst_2.INIT_RAM_25 = 256'h00000810010000400100040808300C30218410081008210410081018200C6020;
defparam prom_inst_2.INIT_RAM_26 = 256'h0180030004300060000000000180031800C00040018018C00380030838C00000;
defparam prom_inst_2.INIT_RAM_27 = 256'h1018000001000100010000000000000000000000000000200180000000C00300;
defparam prom_inst_2.INIT_RAM_28 = 256'h1008200C101828341020061014081408200C0910301810204020300830080240;
defparam prom_inst_2.INIT_RAM_29 = 256'h10088044200400082004002121042104100810080C301D3810102104200C6020;
defparam prom_inst_2.INIT_RAM_2A = 256'h0000018000000000000000000000000003840000018000000000000001840180;
defparam prom_inst_2.INIT_RAM_2B = 256'h00000C0001800000000000000000000000000000000005200000000003800300;
defparam prom_inst_2.INIT_RAM_2C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_2.INIT_RAM_2D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_2.INIT_RAM_2E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_2.INIT_RAM_2F = 256'h018001800180000001800180018000000000018000001018101810180000FFFF;
defparam prom_inst_2.INIT_RAM_30 = 256'h00FFFF0000F00F00006006000060060018FFC60018FFC6000110FFFF80010000;
defparam prom_inst_2.INIT_RAM_31 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_2.INIT_RAM_32 = 256'h02000000000001800100018000C0020001800020011000100440184001801018;
defparam prom_inst_2.INIT_RAM_33 = 256'h1000018000000380018001803010181008000010001004401800100001001008;
defparam prom_inst_2.INIT_RAM_34 = 256'h200430482C240020031808000100101800044010101860102004100802300E08;
defparam prom_inst_2.INIT_RAM_35 = 256'h0000181801000040010004080420042021841008100821040008301820044020;
defparam prom_inst_2.INIT_RAM_36 = 256'h07E007DC0F7B8060707E3F00000007D873F01FF807E019F02FE00FC819F00000;
defparam prom_inst_2.INIT_RAM_37 = 256'h101800000100010001001FF8783C3C3C781E7C3E1E1E1FFC17E03C787BF00FCE;
defparam prom_inst_2.INIT_RAM_38 = 256'h1008200410182C24102002101608160820040910101810204020100810080460;
defparam prom_inst_2.INIT_RAM_39 = 256'h10088044200400082004002121042104100810080420310C1810210420044020;
defparam prom_inst_2.INIT_RAM_3A = 256'h3FFC07E03C3CF00E7FF8387C703E703E0FE863C607E07FF83FFC07FC0FE407F0;
defparam prom_inst_2.INIT_RAM_3B = 256'h3FE01F3E07F4007CF81F01FEF3CEF3CE7E3E3C3E3C3C1FF0F83E3FFC2FE00FCE;
defparam prom_inst_2.INIT_RAM_3C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_2.INIT_RAM_3D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_2.INIT_RAM_3F = 256'h018001800180000001800180018000000000018000001018101810180000FFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h00FFFF0000E00700004182000040020018FFC60018FFC60000E0FFFF80010000;
defparam prom_inst_3.INIT_RAM_01 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_3.INIT_RAM_02 = 256'h02000000000001800100018000C002000180002020E000103FF810C001801018;
defparam prom_inst_3.INIT_RAM_03 = 256'h10000300000000C003C003C0301008100C00001007D004600C00080001001008;
defparam prom_inst_3.INIT_RAM_04 = 256'h6004304824240020011808000100101800040210011840100004100802100F08;
defparam prom_inst_3.INIT_RAM_05 = 256'h00001008010000C0010002000460064021841018100821040008101860044020;
defparam prom_inst_3.INIT_RAM_06 = 256'h0C300C7C114F0060787E3F0000000C7876181FF00C301B18383018681B180000;
defparam prom_inst_3.INIT_RAM_07 = 256'h101800000100010001001FF8F0383C3C781E7C3E1C1C0FFC1C3066783E18186E;
defparam prom_inst_3.INIT_RAM_08 = 256'h1008600410182424102003101208120830040D20011810204020100800080420;
defparam prom_inst_3.INIT_RAM_09 = 256'h1008804420000008200400212104210410081008064021040830210400044020;
defparam prom_inst_3.INIT_RAM_0A = 256'h3FFC0C30383C700E3FF0387C783E783E1838738E0C303FF03FF80FFC1C340C38;
defparam prom_inst_3.INIT_RAM_0B = 256'h3FF0319C0C3C0038F80E01FE719E719E3C3C1C1C3C3C1198701E3FFC3830186E;
defparam prom_inst_3.INIT_RAM_0C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_3.INIT_RAM_0D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_3.INIT_RAM_0E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_3.INIT_RAM_0F = 256'h018001800180000001800180018000000000018000001018101810180000FFFF;
defparam prom_inst_3.INIT_RAM_10 = 256'h00FFFF0000E0070000C1830000C00300080C0400080004000000FFFF80010000;
defparam prom_inst_3.INIT_RAM_11 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_3.INIT_RAM_12 = 256'h0100000000000180010002C000C0030001800060180000600640000001801018;
defparam prom_inst_3.INIT_RAM_13 = 256'h180006007FFE006003C003C030100C30040007100C7004200780080001001008;
defparam prom_inst_3.INIT_RAM_14 = 256'h400430C824640020009808000100101800040610031840100004100802100988;
defparam prom_inst_3.INIT_RAM_15 = 256'h0000000001000080010003000240024023841810100801000010101840042020;
defparam prom_inst_3.INIT_RAM_16 = 256'h1818183811C600600C180E00018018381C08004018181C0C301010381C0C0000;
defparam prom_inst_3.INIT_RAM_17 = 256'h101800200100010001000818201818102004100810180020181843401C041038;
defparam prom_inst_3.INIT_RAM_18 = 256'h1008400410182464102001101208120810000520031810204020100800080420;
defparam prom_inst_3.INIT_RAM_19 = 256'h1008804420000008200400212104210410081008024061040820010000042020;
defparam prom_inst_3.INIT_RAM_1A = 256'h1018181810183814102024101C081C083018511A1818102020601810101C0800;
defparam prom_inst_3.INIT_RAM_1B = 256'h1810608C180C00102004004221042104100808081810310C2008210430101038;
defparam prom_inst_3.INIT_RAM_1C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_3.INIT_RAM_1D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_3.INIT_RAM_1E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_3.INIT_RAM_1F = 256'h018001800180000001800180018000000000018000001018101810180000FFFF;
defparam prom_inst_3.INIT_RAM_20 = 256'h7DFFFFBE7DE007BE00818100008001000C0C0C000C000C000000FFFF80010000;
defparam prom_inst_3.INIT_RAM_21 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_3.INIT_RAM_22 = 256'h0100000000000100010002400080030001000040060003C00240000001801018;
defparam prom_inst_3.INIT_RAM_23 = 256'h08001C000000003803C003C0283007E004000FD0181004200780040001001008;
defparam prom_inst_3.INIT_RAM_24 = 256'h400630882644002000D8080001001018000406100318401000040C0802100888;
defparam prom_inst_3.INIT_RAM_25 = 256'h00000000010000800100010002C0038022440810100801000030181840062020;
defparam prom_inst_3.INIT_RAM_26 = 256'h100810181082006006180C0001801018180C0040100C1C04300830181C040000;
defparam prom_inst_3.INIT_RAM_27 = 256'h101800F00100010001000C1820100C302004100810180020100801C01C062018;
defparam prom_inst_3.INIT_RAM_28 = 256'h1008400610182644102001D0110811080C0007600318102000200C0800080420;
defparam prom_inst_3.INIT_RAM_29 = 256'h1010804460000008200400202104210410081008038041060460010000042020;
defparam prom_inst_3.INIT_RAM_2A = 256'h1018100810182814102026101408140820084912100C102020601010300C0800;
defparam prom_inst_3.INIT_RAM_2B = 256'h1810408C100C00102004004221042104100808080C3021041008210430082018;
defparam prom_inst_3.INIT_RAM_2C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_3.INIT_RAM_2D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_3.INIT_RAM_2E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_3.INIT_RAM_2F = 256'h018001800180000001800180018000000000018000001018101810180000FFFF;
defparam prom_inst_3.INIT_RAM_30 = 256'hFFFFFFFFFFC003FF0F8FF1F00F8FF1F00C0C0C000C000C000000FFFF80010000;
defparam prom_inst_3.INIT_RAM_31 = 256'h1FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF8;
defparam prom_inst_3.INIT_RAM_32 = 256'h010000003FFC00003FFC0460008003000000004001800E000240000001801FF8;
defparam prom_inst_3.INIT_RAM_33 = 256'h060030000000000C018001802C2007E004001850100004100C00060001001008;
defparam prom_inst_3.INIT_RAM_34 = 256'h400231882244002001F8080001001FF8000407F003F84010000407F804180888;
defparam prom_inst_3.INIT_RAM_35 = 256'h00000000010001800100018001800180224408101008010003E00E1840023020;
defparam prom_inst_3.INIT_RAM_36 = 256'h200C10181082006003180C000180101818040040300418022008201818020000;
defparam prom_inst_3.INIT_RAM_37 = 256'h1FF83098010001000180060810100460218C181010180020101800C018022008;
defparam prom_inst_3.INIT_RAM_38 = 256'h100840021FF82244102001F01108110807E007E003F81020002007F80FF80830;
defparam prom_inst_3.INIT_RAM_39 = 256'h1070807C7FC00FF820FC1FE02104210418081008018041020440010000043020;
defparam prom_inst_3.INIT_RAM_3A = 256'h1018200C101828141020221016081608200809103004102020601010200C0800;
defparam prom_inst_3.INIT_RAM_3B = 256'h1810404C10040010200400422104210410080808046021041010210420082008;
defparam prom_inst_3.INIT_RAM_3C = 256'h0003C0001FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF8;
defparam prom_inst_3.INIT_RAM_3D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_3.INIT_RAM_3E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFF01FFFF80FFFFFFFF01FFFF80FF8001FF0180FFFF1FF81FF81FF80000FFFF;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFC003FF0F8FF1F00F8FF1F0040C0800040008000000FFFF80010000;
defparam prom_inst_4.INIT_RAM_01 = 256'h1FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF8;
defparam prom_inst_4.INIT_RAM_02 = 256'h008000003FFC00003FFC042000800300000000E0007018000240000001801FF8;
defparam prom_inst_4.INIT_RAM_03 = 256'h030070000000000E0000000026E00C3006001070100004100800030001001008;
defparam prom_inst_4.INIT_RAM_04 = 256'h4002310822C400200338080001001FF8000407F003F8401000041FF804080888;
defparam prom_inst_4.INIT_RAM_05 = 256'h00000000010001000100008001800180224C0830100801000F0003F840021C20;
defparam prom_inst_4.INIT_RAM_06 = 256'h200410181082006001980C00018010181004004020041802200C200818020000;
defparam prom_inst_4.INIT_RAM_07 = 256'h1FF8110801000100008002001030024031880810101800200010004018022008;
defparam prom_inst_4.INIT_RAM_08 = 256'h100840021FF822C410200310118811880FE00D2003F8102000201FF81FF80810;
defparam prom_inst_4.INIT_RAM_09 = 256'h1FC0807C7FC01FF823FC3FE0210421041C081008018041020640010000041C20;
defparam prom_inst_4.INIT_RAM_0A = 256'h1018200410182C24102003101208120830040520200410202060181020040800;
defparam prom_inst_4.INIT_RAM_0B = 256'h1810C04C200400102004004221042104100808080240210418102104200C2008;
defparam prom_inst_4.INIT_RAM_0C = 256'h0003C0001FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF81FF8;
defparam prom_inst_4.INIT_RAM_0D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_4.INIT_RAM_0E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_4.INIT_RAM_0F = 256'hFFFF01FFFF80FFFFFFFF01FFFF80FF8001FF0180FFFF1FF81FF81FF80000FFFF;
defparam prom_inst_4.INIT_RAM_10 = 256'h7DFFFFBE7DE007BE008181000080010006001800060018000000FFFF80010000;
defparam prom_inst_4.INIT_RAM_11 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_4.INIT_RAM_12 = 256'h00800000000000000100000000800300000010B0001810000240000001001018;
defparam prom_inst_4.INIT_RAM_13 = 256'h01001800000000180000000023C0181002003030100004181000010001001008;
defparam prom_inst_4.INIT_RAM_14 = 256'h400631082284002006180804010010187E040610031840100004300804080888;
defparam prom_inst_4.INIT_RAM_15 = 256'h0000000001000100010000C001000380224C0C20100801001800031840060FE0;
defparam prom_inst_4.INIT_RAM_16 = 256'h200410181082006000D80C000180101810040040200418020004600818020000;
defparam prom_inst_4.INIT_RAM_17 = 256'h10181F040600010000E0030018200380118808101018002000F0004018026008;
defparam prom_inst_4.INIT_RAM_18 = 256'h1008400610182284102002101088108818000930031810200020300830080810;
defparam prom_inst_4.INIT_RAM_19 = 256'h10C08044600030082204602021042104161810080380410602C0010000040FE0;
defparam prom_inst_4.INIT_RAM_1A = 256'h101820041018242410200190130813081C0007602004102020600FF060040FE0;
defparam prom_inst_4.INIT_RAM_1B = 256'h1810804C20000010200400402104210410080808038061040830210400046008;
defparam prom_inst_4.INIT_RAM_1C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_4.INIT_RAM_1D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_4.INIT_RAM_1E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_4.INIT_RAM_1F = 256'h018001800180018000000000000001800180018000001018101810180000FFFF;
defparam prom_inst_4.INIT_RAM_20 = 256'h01FFFF8001E0078000C1830000C0030003001000030010000000FFFF80010000;
defparam prom_inst_4.INIT_RAM_21 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_4.INIT_RAM_22 = 256'h00800000000000000100000000800300000019900F0410001FF8000001001018;
defparam prom_inst_4.INIT_RAM_23 = 256'h01000C007FFE0070000000002000101802002030100004081000018001001008;
defparam prom_inst_4.INIT_RAM_24 = 256'h400632082184402004180804010010187F04061003184010000420080FF80888;
defparam prom_inst_4.INIT_RAM_25 = 256'h0000000001000300010000400100024026480420100801001000061840060020;
defparam prom_inst_4.INIT_RAM_26 = 256'h200410181082006000380C0001801018100400403FFC18020004400818020000;
defparam prom_inst_4.INIT_RAM_27 = 256'h10180E000700010000C0010008200180138808201018002007C0004018024008;
defparam prom_inst_4.INIT_RAM_28 = 256'h10084006101821841020061010C810C830000910031810200020200820081FF0;
defparam prom_inst_4.INIT_RAM_29 = 256'h1060804460002008260440202104210413F01008024061040280010000040020;
defparam prom_inst_4.INIT_RAM_2A = 256'h101820041FF82424102001F01108110807E007E03FFC102020600FF060040FF0;
defparam prom_inst_4.INIT_RAM_2B = 256'h1830807C3FC007F021FC3FC02104210418080808018061040820210400044008;
defparam prom_inst_4.INIT_RAM_2C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_4.INIT_RAM_2D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_4.INIT_RAM_2E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_4.INIT_RAM_2F = 256'h018001800180018000000000000001800180018000001018101810180000FFFF;
defparam prom_inst_4.INIT_RAM_30 = 256'h00FFFF0000E00700004182000040020001807800018078000000FFFF80010000;
defparam prom_inst_4.INIT_RAM_31 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_4.INIT_RAM_32 = 256'h0040000000000000010000000080030000000910088010081FFC000000001018;
defparam prom_inst_4.INIT_RAM_33 = 256'h010007007FFC00C000000000100010080200201030001FF8100000C001001008;
defparam prom_inst_4.INIT_RAM_34 = 256'h60043208218440200C180804010010182004001000184010000460080FFC0988;
defparam prom_inst_4.INIT_RAM_35 = 256'h00000000010002000100106001000660346804201008010030000C1860040020;
defparam prom_inst_4.INIT_RAM_36 = 256'h200410181082006000780C000180101810040040000418020004400818020000;
defparam prom_inst_4.INIT_RAM_37 = 256'h1018000001000100008000800840038012C80420101800200C00004018026008;
defparam prom_inst_4.INIT_RAM_38 = 256'h1008600410182184102004101048104820001118001810200020600860081FF8;
defparam prom_inst_4.INIT_RAM_39 = 256'h10308044200060082404C0202104210410E01008066021040180010000040020;
defparam prom_inst_4.INIT_RAM_3A = 256'h101820041018264410200310108810881F000D20000410202060181060040818;
defparam prom_inst_4.INIT_RAM_3B = 256'h1FE0804C3FC00C1023847040210421041E180808038061040420010000046008;
defparam prom_inst_4.INIT_RAM_3C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_4.INIT_RAM_3D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_4.INIT_RAM_3E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_4.INIT_RAM_3F = 256'h018001800180018000000000000001800180018000001018101810180000FFFF;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h00FFFF0000F00F00006006000060060000E1DE0000E1DE000000FFFF80010000;
defparam prom_inst_5.INIT_RAM_01 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_5.INIT_RAM_02 = 256'h0040000000000000010000000080030000000B18108010080260000000001018;
defparam prom_inst_5.INIT_RAM_03 = 256'h0000018000000180000000001000100802002010100004003000004001001008;
defparam prom_inst_5.INIT_RAM_04 = 256'h2004360820044020081808040100101820040010201840100004400808041F08;
defparam prom_inst_5.INIT_RAM_05 = 256'h0000000001000200010010200100042014280440100801002000081820040020;
defparam prom_inst_5.INIT_RAM_06 = 256'h200410181082006000D80C000180101810040040000418020004600818020000;
defparam prom_inst_5.INIT_RAM_07 = 256'h1018000001000100010000C00C40024012480420101800201000004018022008;
defparam prom_inst_5.INIT_RAM_08 = 256'h100820041018200410200C101048104820001108201810200020400840081008;
defparam prom_inst_5.INIT_RAM_09 = 256'h10108044200040082404802021042104100010080420310C0180010000040020;
defparam prom_inst_5.INIT_RAM_0A = 256'h10182004101822441020021010C810C83000091000041020006030106004080C;
defparam prom_inst_5.INIT_RAM_0B = 256'h1FC0804C20001010220440402104210417F00808024061040460010000042008;
defparam prom_inst_5.INIT_RAM_0C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_5.INIT_RAM_0D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_5.INIT_RAM_0E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_5.INIT_RAM_0F = 256'h018001800180018000000000000001800180018000001018101810180000FFFF;
defparam prom_inst_5.INIT_RAM_10 = 256'h007FFE00007E7E0000300C0000300C00007F8F00007F8F000000FFFF80010000;
defparam prom_inst_5.INIT_RAM_11 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_5.INIT_RAM_12 = 256'h0040000000000000010000000080030000000A08104018180260000000001018;
defparam prom_inst_5.INIT_RAM_13 = 256'h000000C00000030001C000001000100803002010100004001000002001001018;
defparam prom_inst_5.INIT_RAM_14 = 256'h200434082004402008180804010010182004001020182010000C400808040008;
defparam prom_inst_5.INIT_RAM_15 = 256'h00000000010006000100103001000C301428024010080100200C181820040020;
defparam prom_inst_5.INIT_RAM_16 = 256'h200410181082006001980C00018010181804004000041802000C200818020000;
defparam prom_inst_5.INIT_RAM_17 = 256'h1018000001000100010000400440066012580460101800201000004018022008;
defparam prom_inst_5.INIT_RAM_18 = 256'h1008200410182004102008101028102820001108201810200020400840081008;
defparam prom_inst_5.INIT_RAM_19 = 256'h10188044200040082404802021042104100010080C30191801800100000C0020;
defparam prom_inst_5.INIT_RAM_1A = 256'h1018200410182244102004101048104820001910000410200060201020040804;
defparam prom_inst_5.INIT_RAM_1B = 256'h1860C04C20001010220440402104210410E008080660210406400100000C2008;
defparam prom_inst_5.INIT_RAM_1C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_5.INIT_RAM_1D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_5.INIT_RAM_1E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_5.INIT_RAM_1F = 256'h018001800180018000000000000001800180018000001018101810180000FFFF;
defparam prom_inst_5.INIT_RAM_20 = 256'h01FFFF8001FFFF80001C3800001C380000000F8000000F800000FFFF80010000;
defparam prom_inst_5.INIT_RAM_21 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_5.INIT_RAM_22 = 256'h00200000000000000100000000C0030000000E18104008180220000000001018;
defparam prom_inst_5.INIT_RAM_23 = 256'h0000006000000E0001C000001800100801003020100004001000003001001810;
defparam prom_inst_5.INIT_RAM_24 = 256'h300C3408200440201818080401001018200C0010201820102008600818040008;
defparam prom_inst_5.INIT_RAM_25 = 256'h000000000100040001001010010008101428024010080100300C1018300C0020;
defparam prom_inst_5.INIT_RAM_26 = 256'h200C10181082006003180C0001801018180C0040000C18020008201818020000;
defparam prom_inst_5.INIT_RAM_27 = 256'h10180000010001000100106004800C301650024010180020100800401C062018;
defparam prom_inst_5.INIT_RAM_28 = 256'h1008300C10182004102108101028102820003108201810300020600860083008;
defparam prom_inst_5.INIT_RAM_29 = 256'h1008C044100460082404C020210421041000100808100FF00084010020080020;
defparam prom_inst_5.INIT_RAM_2A = 256'h1018200C1018228410200C101068106820001108000C102000602010200C0804;
defparam prom_inst_5.INIT_RAM_2B = 256'h1830404C300010102604404021042104100008080C30210402C0010000082018;
defparam prom_inst_5.INIT_RAM_2C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_5.INIT_RAM_2D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_5.INIT_RAM_2E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_5.INIT_RAM_2F = 256'h018001800180018000000000000001800180018000001018101810180000FFFF;
defparam prom_inst_5.INIT_RAM_30 = 256'h03DFFBC003DFFBC0C007E003C007E00300000FC000000FC00000FFFF80010000;
defparam prom_inst_5.INIT_RAM_31 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_5.INIT_RAM_32 = 256'h002003C0000000000100000000C002000000041010400FE80220000000001018;
defparam prom_inst_5.INIT_RAM_33 = 256'h000000380000180000E003C00C00181801001020180804001000001801000810;
defparam prom_inst_5.INIT_RAM_34 = 256'h1008380820044020101808040100101820080010201830106018200810020008;
defparam prom_inst_5.INIT_RAM_35 = 256'h00000000010004000100101801001018182802C010180100100C301810080020;
defparam prom_inst_5.INIT_RAM_36 = 256'h100810181082006006180C00018010181C08004000081C04200830181C040000;
defparam prom_inst_5.INIT_RAM_37 = 256'h101800000100010001001030068008100C70024018180020100800401C0C1038;
defparam prom_inst_5.INIT_RAM_38 = 256'h1008100810182004102318101038103820022104201810100020200820082004;
defparam prom_inst_5.INIT_RAM_39 = 256'h100840C410042008240440202104210410001008101807C00084010060180020;
defparam prom_inst_5.INIT_RAM_3A = 256'h1018100810182184102208101028102820001108000810200060201030080804;
defparam prom_inst_5.INIT_RAM_3B = 256'h1810408C10041010220440402104210410000808081021040280010020081038;
defparam prom_inst_5.INIT_RAM_3C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_5.INIT_RAM_3D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F001F000F0007000300010000;
defparam prom_inst_5.INIT_RAM_3E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_5.INIT_RAM_3F = 256'h018001800180018000000000000001800180018000001018101810180000FFFF;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h07C7E3E007C7E3E0C0018003C0018003000007E0000007E00000FFFF80010000;
defparam prom_inst_6.INIT_RAM_01 = 256'h1018101810181018101810181018101810181018101810181018101810181018;
defparam prom_inst_6.INIT_RAM_02 = 256'h002003C0000000000100000000C0020000000610108003C80220000001801018;
defparam prom_inst_6.INIT_RAM_03 = 256'h03C0000C0000300000E003C00400081001001060081804000808100C01000C30;
defparam prom_inst_6.INIT_RAM_04 = 256'h181838082004402010180C080100101820180010201818103010300810020010;
defparam prom_inst_6.INIT_RAM_05 = 256'h0000000001000C0001001008010030081838038008100100101C201818180020;
defparam prom_inst_6.INIT_RAM_06 = 256'h18181018108200600C180C00018010181610004020181C0C301010381C0C0000;
defparam prom_inst_6.INIT_RAM_07 = 256'h101800000100010001001010028010180C3002C01C102020100800401E181868;
defparam prom_inst_6.INIT_RAM_08 = 256'h10081818101820041023101010181018300C2104201810180020300830082004;
defparam prom_inst_6.INIT_RAM_09 = 256'h10044084080C30082204602021042104100010083008010000C4010030100020;
defparam prom_inst_6.INIT_RAM_0A = 256'h101818181018218410221810103810382004210C201810100060301010180C04;
defparam prom_inst_6.INIT_RAM_0B = 256'h1818608C180C18102204404021042104100008081018310C0380010030101868;
defparam prom_inst_6.INIT_RAM_0C = 256'h0003C00010181018101810181018101810181018101810181018101810181018;
defparam prom_inst_6.INIT_RAM_0D = 256'h7FFF3FFF1FFF0FFF07FF03FF01FF00FF007F003F003F001F0007000300010000;
defparam prom_inst_6.INIT_RAM_0E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_6.INIT_RAM_0F = 256'h018001800180018000000000000001800180018000001018101810180000FFFF;
defparam prom_inst_6.INIT_RAM_10 = 256'h0F8181F00F8181F0C0018003C0018003000003F0000003F00000FFFF80010000;
defparam prom_inst_6.INIT_RAM_11 = 256'h7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C;
defparam prom_inst_6.INIT_RAM_12 = 256'h001003C000000000010000000040060000001A30188001000220000003C07C3C;
defparam prom_inst_6.INIT_RAM_13 = 256'h03C000040000200000E003C003100C20018008C00C301F000C381FFC1FF80460;
defparam prom_inst_6.INIT_RAM_14 = 256'h0C30383CF81E7FFC707C06381FF87C3C307003FC3FFC0FFC18601FFC7C0F0010;
defparam prom_inst_6.INIT_RAM_15 = 256'h000000000100080001001FF80FF0783E181801800C300FF00C3CE07C0C3003F8;
defparam prom_inst_6.INIT_RAM_16 = 256'h0C30383C71870FF8787C0C000FF0383C93F01FF838303B181830186E3B180000;
defparam prom_inst_6.INIT_RAM_17 = 256'h7C3C00000100010001001FF803007C3C0C3003803630306018380FF81BF00FC8;
defparam prom_inst_6.INIT_RAM_18 = 256'h3C3C0C307C3CF81E7C13707C7C1E7C1E181CE3C73FFC7FFE01FC1FFC1FFCF81E;
defparam prom_inst_6.INIT_RAM_19 = 256'h7E06618E0C181FFCFBFF3FF0FFFEFFFE3F007FFC783E03C000440FF0186003F8;
defparam prom_inst_6.INIT_RAM_1A = 256'h3C3C0C303C3C783E7C32707C7C1E7C1E381C63C638307FFE01FC1FFC1C303F08;
defparam prom_inst_6.INIT_RAM_1B = 256'h3E0C319E0C180FF8FBFE7FE0FFFE7FFE3F007FFE7C3C119801800FF018300FC8;
defparam prom_inst_6.INIT_RAM_1C = 256'h0003C0007C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C7C3C;
defparam prom_inst_6.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_6.INIT_RAM_1F = 256'h018001800180018000000000000001800180018000007C3C7C3C7C3C0000FFFF;
defparam prom_inst_6.INIT_RAM_20 = 256'h1F03C0F81F03C0F8C0018003C0018003000001F8000001F80000FFFF80010000;
defparam prom_inst_6.INIT_RAM_21 = 256'h7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E;
defparam prom_inst_6.INIT_RAM_22 = 256'h001003C000000000000000000060060000001BE00F0001000220000003807C7E;
defparam prom_inst_6.INIT_RAM_23 = 256'h03C0000000000000006003C001F007E000800F8007E01F8007E01FFC1FF807C0;
defparam prom_inst_6.INIT_RAM_24 = 256'h07E0307EFC3F7FFC707E03F01FF87C7E1FE003FC3FFE07FC0FC00FFE7E1F8830;
defparam prom_inst_6.INIT_RAM_25 = 256'h000000000100080001001FF80FF07C3E1818018007E00FF007E4C07E07E003FC;
defparam prom_inst_6.INIT_RAM_26 = 256'h07E07C7E718F8FF8707E0C080FF07C7E90C01FF80FE079F00FE00FCE79F00000;
defparam prom_inst_6.INIT_RAM_27 = 256'h7C7E00000100010001001FF803007C3E0C30018073E01FC00FE80FFC18C00308;
defparam prom_inst_6.INIT_RAM_28 = 256'h7C7E07E07C7EFC3F7C1FF07CFC0EFC0E0FF0C3C73FFE7FFE03FC0FFE0FFEFC3F;
defparam prom_inst_6.INIT_RAM_29 = 256'h7E073F1F07F00FFEF9FF1FF0FFFFFFFF7F807FFE7C3E07E0003C0FF00FC003FC;
defparam prom_inst_6.INIT_RAM_2A = 256'h7C7E07E07C7EFC3F7C1E707C7C0E7C0E1FF8E3C70FE07FFE03FC0FFC0FE079F8;
defparam prom_inst_6.INIT_RAM_2B = 256'h3E0C1F3F07F007FCF9FF1FE0FFFFFFFF7F007FFE7C3E1FF001000FF00FE00308;
defparam prom_inst_6.INIT_RAM_2C = 256'h0003C0007C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E7C7E;
defparam prom_inst_6.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_2E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C0008000FFFF;
defparam prom_inst_6.INIT_RAM_2F = 256'h018001800180018000000000000001800180018000007C7E7C7E7C7E0000FFFF;
defparam prom_inst_6.INIT_RAM_30 = 256'h3E03C07C3E03C07C6001800660018006000000FC000000FC0000FFFF80010000;
defparam prom_inst_6.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_32 = 256'h0010018000000000000000000060040000000080000001000220000001800000;
defparam prom_inst_6.INIT_RAM_33 = 256'h0180000000000000006001800060018000000200018000000180000000000180;
defparam prom_inst_6.INIT_RAM_34 = 256'h0180000000000000000000C00000000003000000000000000300000000000C60;
defparam prom_inst_6.INIT_RAM_35 = 256'h0000000001001800010000000000000000000000018000000180000001800000;
defparam prom_inst_6.INIT_RAM_36 = 256'h0180000000000000000006080000000010000000038000C00380030000C00000;
defparam prom_inst_6.INIT_RAM_37 = 256'h000000000100010001000000010000000000000000C003000180000018000008;
defparam prom_inst_6.INIT_RAM_38 = 256'h0000018000000000000400000000000003800000000040020000000000000000;
defparam prom_inst_6.INIT_RAM_39 = 256'h00000C0001C00000000000008000000000004000000000000018000003000000;
defparam prom_inst_6.INIT_RAM_3A = 256'h0000018000000000000C00000000000003800000038040020000000001800060;
defparam prom_inst_6.INIT_RAM_3B = 256'h00000C0001800000000000008000000000004000000003200084000003800008;
defparam prom_inst_6.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3E = 256'hFFFEFFFCFFF8FFF0FFE0FFC0FF80FF00FE00FC00F800F000E000C00080000000;
defparam prom_inst_6.INIT_RAM_3F = 256'h018001800180018000000000000001800180018000000000000000000000FFFF;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h3C03C03C3C03C03C600000066000000600000078000000780000FFFF80010000;
defparam prom_inst_7.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_02 = 256'h00080000000000000000000000200C0000000000000001000220000000000000;
defparam prom_inst_7.INIT_RAM_03 = 256'h0000000000000000003000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_04 = 256'h00000000000000000000000000000000000000000000000000000000000007C0;
defparam prom_inst_7.INIT_RAM_05 = 256'h0000000001001000010000000000000000000000000000000000000000400000;
defparam prom_inst_7.INIT_RAM_06 = 256'h0000000000000000000006180000000010000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_07 = 256'h0000000001800100010000000100000000000000000000000000000018000008;
defparam prom_inst_7.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000040020000000000000000;
defparam prom_inst_7.INIT_RAM_09 = 256'h0000000000000000000000008000000000004000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000040020000000000000000;
defparam prom_inst_7.INIT_RAM_0B = 256'h0000000000000000000000008000000000004000000001000084000000000008;
defparam prom_inst_7.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0F = 256'h0180018001800180000000000000018001800180000000000000000000000000;
defparam prom_inst_7.INIT_RAM_10 = 256'h1803C0181803C0183800001C3800001C00000030000000300000FFFF80010000;
defparam prom_inst_7.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_12 = 256'h0008000000000000000000000030080000000000000001000000000000000000;
defparam prom_inst_7.INIT_RAM_13 = 256'h0000000000000000003000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_15 = 256'h0000000001001000010000000000000000000000000000000000000067E00000;
defparam prom_inst_7.INIT_RAM_16 = 256'h0000000000000000000006300000000010000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_17 = 256'h0000000000800100010000000080000000000000000000000000000018000008;
defparam prom_inst_7.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000040020000000000000000;
defparam prom_inst_7.INIT_RAM_19 = 256'h0000000000000000000000008000000000004000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000040020000000000000000;
defparam prom_inst_7.INIT_RAM_1B = 256'h00000000000000000000000080000000000040000000010000C4000000000008;
defparam prom_inst_7.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1F = 256'h0180018001800180000000000000018001800180000000000000000000000000;
defparam prom_inst_7.INIT_RAM_20 = 256'h0003C0000003C0001F8001F81F8001F800000000000000000000FFFF80010000;
defparam prom_inst_7.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_22 = 256'h0000000000000000000000000010080000000000000000800000000000000000;
defparam prom_inst_7.INIT_RAM_23 = 256'h0000000000000000001000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_25 = 256'h0000000001F000000F000000000000000000000000000000000000003EF00000;
defparam prom_inst_7.INIT_RAM_26 = 256'h0000000000000000000003E00000000018000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_27 = 256'h0000000000E00100070000000080000000000000000000000000000018000008;
defparam prom_inst_7.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000040020000000000000000;
defparam prom_inst_7.INIT_RAM_29 = 256'h0000000000000000000000008000000000004000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000040020000000000000000;
defparam prom_inst_7.INIT_RAM_2B = 256'h0000000000000000000000008000000000004000000001000044000000000008;
defparam prom_inst_7.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2F = 256'h0180018001800180000000000000018001800180000000000000000000000000;
defparam prom_inst_7.INIT_RAM_30 = 256'h0001800000018000078001E0078001E000000000000000000000FFFFFFFF0000;
defparam prom_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000010080000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_35 = 256'h0000000001F000000F0000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_36 = 256'h0000000000000000000001C00000000008000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_37 = 256'h0000000000600100060000000080000000000000000000000000000018000008;
defparam prom_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000040020000000000000000;
defparam prom_inst_7.INIT_RAM_39 = 256'h0000000000000000000000008000000000004000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3B = 256'h000000000000000000000000000000000000000000000FE0007C000000000008;
defparam prom_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3F = 256'h0180018001800180000000000000018001800180000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(prom_inst_4_dout[0]),
  .I1(prom_inst_5_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(prom_inst_6_dout[0]),
  .I1(prom_inst_7_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_1)
);
MUX2 mux_inst_6 (
  .O(dout[0]),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_0)
);
endmodule //table_FONT
