//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-3
//Part Number: GW2AR-LV18EQ144C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Fri Nov 10 08:56:16 2023

module bme240_i2cmem (dout, clk, oce, ce, reset, ad);

output [8:0] dout;
input clk;
input oce;
input ce;
input reset;
input [8:0] ad;

wire [26:0] promx9_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROMX9 promx9_inst_0 (
    .DO({promx9_inst_0_dout_w[26:0],dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,gw_gnd,ad[8:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_0.READ_MODE = 1'b0;
defparam promx9_inst_0.BIT_WIDTH = 9;
defparam promx9_inst_0.RESET_MODE = "SYNC";
defparam promx9_inst_0.INIT_RAM_00 = 288'h287D3E4105BBD1DDF100063E9F202BC9DDF10000001F4F9840C1F5F97C1DFF1F9341DDF1;
defparam promx9_inst_0.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_02 = 288'h00000A1F4F9A0009F5F97C1DFF1F93CDDDF1000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_04 = 288'hF97C1DFF1F93E9DDF1F97C1DFF1F93E5DDF1F97C1DFF1F93E1DDF1F97C1DFF1F93DDDDF1;
defparam promx9_inst_0.INIT_RAM_05 = 288'hF97C1DFF1F93F9DDF1F97C1DFF1F93F5DDF1F97C1DFF1F93F1DDF1F97C1DFF1F93EDDDF1;
defparam promx9_inst_0.INIT_RAM_06 = 288'h00000000000000000000000000000000000000000000000000000000000000000001E1F4;
defparam promx9_inst_0.INIT_RAM_07 = 288'hF97C1DFF1F9225DDF1F97C1DFF1F9221DDF1000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_08 = 288'hF97C1DFF1F9235DDF1F97C1DFF1F9231DDF1F97C1DFF1F922DDDF1F97C1DFF1F9229DDF1;
defparam promx9_inst_0.INIT_RAM_09 = 288'hF97C1DFF1F9245DDF1F97C1DFF1F9241DDF1F97C1DFF1F923DDDF1F97C1DFF1F9239DDF1;
defparam promx9_inst_0.INIT_RAM_0A = 288'hF97C1DFF1F9255DDF1F97C1DFF1F9251DDF1F97C1DFF1F924DDDF1F97C1DFF1F9249DDF1;
defparam promx9_inst_0.INIT_RAM_0B = 288'hF97C1DFF1F9265DDF1F97C1DFF1F9261DDF1F97C1DFF1F925DDDF1F97C1DFF1F9259DDF1;
defparam promx9_inst_0.INIT_RAM_0C = 288'hF97C1DFF1F9275DDF1F97C1DFF1F9271DDF1F97C1DFF1F926DDDF1F97C1DFF1F9269DDF1;
defparam promx9_inst_0.INIT_RAM_0D = 288'hF97C1DFF1F9385DDF1F97C1DFF1F9285DDF1F97C1DFF1F927DDDF1F97C1DFF1F9279DDF1;
defparam promx9_inst_0.INIT_RAM_0E = 288'hF97C1DFF1F9395DDF1F97C1DFF1F9391DDF1F97C1DFF1F938DDDF1F97C1DFF1F9389DDF1;
defparam promx9_inst_0.INIT_RAM_0F = 288'h0000000000000000000000000000000001F4F97C1DFF1F939DDDF1F97C1DFF1F9399DDF1;

endmodule //bme240_i2cmem
