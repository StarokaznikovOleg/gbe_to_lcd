//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2AR-LV18EQ144C8/I7
//Device: GW2AR-18C
//Created Time: Fri Nov 04 21:15:09 2022

module logo_rom (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [16:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [0:0] prom_inst_4_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire mux_o_0;
wire mux_o_1;
wire mux_o_3;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_0.INIT = 16'h0002;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_1.INIT = 16'h0008;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_2.INIT = 16'h0020;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_3.INIT = 16'h0080;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_4.INIT = 16'h0200;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000003E00000000000000000000000000000000000078000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000003C0000000000000000000000000000000000007C000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000007C0000000000000000000000000000000000003E000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000007C0000000000000000000000000000000000003E000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h000000000001F80000000000000000000000000000000000001F800000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h000000000003F80000000000000000000000000000000000001FC00000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h000000000003F00000000000000000000000000000000000000FC00000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h000000000007E00000000000000000000000000000000000000FE00000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h00000000000FE007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE007F00000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'h00000000001FC007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE003F80000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h00000000003F800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001F80000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h00000000003F800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001F80000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h00000000007F800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FC0000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h00000000007E003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC007E0000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000000FC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003F0000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000000001F8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001F8000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000003F8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FC000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h000000000FF000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FF000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h000000003FE001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007F800000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h000000007FC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FE00000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h00000000FF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001FF00000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h00000003FF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFC0000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000FFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FE0000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h0000003FF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFC000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h000000FFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FF000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h000000FFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FF000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h000007FF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFC00000;
defparam prom_inst_0.INIT_RAM_24 = 256'h00001FFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFF80000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0001FFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFF8000;
defparam prom_inst_0.INIT_RAM_26 = 256'h001FFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFF000;
defparam prom_inst_0.INIT_RAM_27 = 256'h01FFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FFFF00;
defparam prom_inst_0.INIT_RAM_28 = 256'h03FFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFC0;
defparam prom_inst_0.INIT_RAM_29 = 256'h0FFFE000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FFC0;
defparam prom_inst_0.INIT_RAM_2A = 256'h0FFC0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000003FF0;
defparam prom_inst_0.INIT_RAM_2B = 256'h0FC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003F0;
defparam prom_inst_0.INIT_RAM_2C = 256'h0FC0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000003F8;
defparam prom_inst_0.INIT_RAM_2D = 256'h0F8000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000003F8;
defparam prom_inst_0.INIT_RAM_2E = 256'h0F8000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000001F0;
defparam prom_inst_0.INIT_RAM_2F = 256'h0F800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00001F0;
defparam prom_inst_0.INIT_RAM_30 = 256'h0F800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00001F0;
defparam prom_inst_0.INIT_RAM_31 = 256'h0F80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001F0;
defparam prom_inst_0.INIT_RAM_32 = 256'h0F8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8001F0;
defparam prom_inst_0.INIT_RAM_33 = 256'h1F803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01F0;
defparam prom_inst_0.INIT_RAM_34 = 256'h1F803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01F0;
defparam prom_inst_0.INIT_RAM_35 = 256'h1F803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01F8;
defparam prom_inst_0.INIT_RAM_36 = 256'h1F807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01F8;
defparam prom_inst_0.INIT_RAM_37 = 256'h1F007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01F8;
defparam prom_inst_0.INIT_RAM_38 = 256'h1F007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00F8;
defparam prom_inst_0.INIT_RAM_39 = 256'h1F007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00F8;
defparam prom_inst_0.INIT_RAM_3A = 256'h1F007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00F8;
defparam prom_inst_0.INIT_RAM_3B = 256'h1F007FFFFFFFC000000000000000000000000000001FFFFFFFFFFFFFFFFE00F8;
defparam prom_inst_0.INIT_RAM_3C = 256'h1F007FFFFFFFC00000000000000000000000000000003FFFFFFFFFFFFFFE00F8;
defparam prom_inst_0.INIT_RAM_3D = 256'h1F007FFFFFFFC00000000000000000000000000000003FFFFFFFFFFFFFFE00F8;
defparam prom_inst_0.INIT_RAM_3E = 256'h1F007FFFFFFFC000000000000000000000000000000007FFFFFFFFFFFFFE00F8;
defparam prom_inst_0.INIT_RAM_3F = 256'h1F007FFFFFFFC000000000000000000000000000000000FFFFFFFFFFFFFE00F8;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h1F01FFFFFFFFC0000000000000000000000000000000003FFFFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_01 = 256'h1F01FFFFFFFFC0000000000000000000000000000000000FFFFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_02 = 256'h1F01FFFFFFFFC00000000000000000000000000000000003FFFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_03 = 256'h1F01FFFFFFFFC00000000000000000000000000000000001FFFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_04 = 256'h1F01FFFFFFFFC00000000000000000000000000000000000FFFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_05 = 256'h1F01FFFFFFFFC000000000000000000000000000000000007FFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_06 = 256'h1F01FFFFFFFFC000000000000000000000000000000000003FFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_07 = 256'h1F01FFFFFFFFC000000000000000000000000000000000003FFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_08 = 256'h1F01FFFFFFFFC000000000000000000000000000000000001FFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_09 = 256'h1F01FFFFFFFFC000000000000000000000000000000000000FFFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_0A = 256'h1F01FFFFFFFFC0000000000000000000000000000000000003FFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_0B = 256'h1F01FFFFFFFFC0000000000000000000000000000000000003FFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_0C = 256'h1F01FFFFFFFFC0000000000000000000000000000000000003FFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_0D = 256'h1F01FFFFFFFFC0000000000000000000000000000000000001FFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_0E = 256'h1F01FFFFFFFFC0000000000000000000000000000000000000FFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_0F = 256'h1F01FFFFFFFFC0000000000000000000000000000000000000FFFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_10 = 256'h1F01FFFFFFFFC00000000000000000000000000000000000007FFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_11 = 256'h1F01FFFFFFFFC00000000000000000000000000000000000007FFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_12 = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFF8001FFFFE000003FFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_13 = 256'h1F01FFFFFFFFFFFFFFFFFF000007FFFFFFFF8001FFFFFE00003FFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_14 = 256'h1F01FFFFFFFFFFFFFFFFFF000007FFFFFFFF8001FFFFFFC0001FFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_15 = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFF8000FFFFFFF8001FFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_16 = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFF8000FFFFFFFC000FFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_17 = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFF8000FFFFFFFE000FFFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_18 = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFFC000FFFFFFFF8007FFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_19 = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFFC000FFFFFFFF8007FFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_1A = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFFC000FFFFFFFFC007FFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_1B = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFFC000FFFFFFFFE003FFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_1C = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFFC000FFFFFFFFE003FFFFFFFF80F8;
defparam prom_inst_1.INIT_RAM_1D = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFFC000FFFFFFFFF003FFFFFFFF80F0;
defparam prom_inst_1.INIT_RAM_1E = 256'h1F01FFFFFFFFFFFFFFFFFF000003FFFFFFFFC000FFFFFFFFFC01FFFFFFFF81F0;
defparam prom_inst_1.INIT_RAM_1F = 256'h0F81FFFFFFFFFFFFFFFFFF800003FFFFFFFFC0007FFFFFFFFE01FFFFFFFF81F0;
defparam prom_inst_1.INIT_RAM_20 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFF007FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_21 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFF007FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_22 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFF807FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_23 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFFC03FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_24 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFFC03FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_25 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFFE03FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_26 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFFE03FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_27 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFFF01FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_28 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0007FFFFFFFFFF01FFFFFFE01F0;
defparam prom_inst_1.INIT_RAM_29 = 256'h0F807FFFFFFFFFFFFFFFFF800001FFFFFFFFC0003FFFFFFFFFFFFFFFFFFE01C0;
defparam prom_inst_1.INIT_RAM_2A = 256'h03C07FFFFFFFFFFFFFFFFF800001FFFFFFFFE0003FFFFFFFFFFFFFFFFFFE03C0;
defparam prom_inst_1.INIT_RAM_2B = 256'h03C07FFFFFFFFFFFFFFFFF800001FFFFFFFFE0003FFFFFFFFFFFFFFFFFFE03C0;
defparam prom_inst_1.INIT_RAM_2C = 256'h03C07FFFFFFFFFFFFFFFFF8000007FFFFFFFE0003FFFFFFFFFFFFFFFFFFC03C0;
defparam prom_inst_1.INIT_RAM_2D = 256'h03C03FFFFFFFFFFFFFFFFF8000007FFFFFFFE0003FFFFFFFFFFFFFFFFFFC03C0;
defparam prom_inst_1.INIT_RAM_2E = 256'h03C03FFFFFFFFFFFFFFFFF8000007FFFFFFFE0003FFFFFFFFFFFFFFFFFFC03C0;
defparam prom_inst_1.INIT_RAM_2F = 256'h03C03FFFFFFFFFFFFFFFFFC000007FFFFFFFE0003FFFFFFFFFFFFFFFFFFC03C0;
defparam prom_inst_1.INIT_RAM_30 = 256'h03C03FFFFFFFFFFFFFFFFFC000007FFFFFFFE0001FFFFFFFFFFFFFFFFFFC03C0;
defparam prom_inst_1.INIT_RAM_31 = 256'h03C03FFFFFFFFFFFFFFFFFC000007FFFFFFFE0001FFFFFFFFFFFFFFFFFFC0380;
defparam prom_inst_1.INIT_RAM_32 = 256'h01E03FFFFFFFFFFFFFFFFFC000007FFFFFFFE0001FFFFFFFFFFFFFFFFFFC0780;
defparam prom_inst_1.INIT_RAM_33 = 256'h01E03FFFFFFFFFFFFFFFFFC000007FFFFFFFE0001FFFFFFFFFFFFFFFFFFC0780;
defparam prom_inst_1.INIT_RAM_34 = 256'h01E03FFFFFFFFFFFFFFFFFC000007FFFFFFFE0001FFFFFFFFFFFFFFFFFFC0780;
defparam prom_inst_1.INIT_RAM_35 = 256'h01E01FFFFFFFFFFFFFFFFFC000007FFFFFFFE0001FFFFFFFFFFFFFFFFFF80780;
defparam prom_inst_1.INIT_RAM_36 = 256'h01E01FFFFFFFFFFFFFFFFFC000007FFFFFFFE0001FFFFFFFFFFFFFFFFFF80780;
defparam prom_inst_1.INIT_RAM_37 = 256'h01E01FFFFFFFFFFFFFFFFFC000003FFFFFFFF0001FFFFFFFFFFFFFFFFFF80780;
defparam prom_inst_1.INIT_RAM_38 = 256'h01E01FFFFFFFFFFFFFFFFFC000003FFFFFFFF0000FFFFFFFFFFFFFFFFFF80700;
defparam prom_inst_1.INIT_RAM_39 = 256'h00F01FFFFFFFFFFFFFFFFFC000003FFFFFFFF0000FFFFFFFFFFFFFFFFFF80F00;
defparam prom_inst_1.INIT_RAM_3A = 256'h00F01FFFFFFFFFFFFFFFFFC000003FFFFFFFF0000FFFFFFFFFFFFFFFFFF80F00;
defparam prom_inst_1.INIT_RAM_3B = 256'h00F01FFFFFFFFFFFFFFFFFC000003FFFFFFFF0000FFFFFFFFFFFFFFFFFF00F00;
defparam prom_inst_1.INIT_RAM_3C = 256'h00F00FFFFFFFFFFFFFFFFFC000003FFFFFFFF0000FFFFFFFFFFFFFFFFFF00F00;
defparam prom_inst_1.INIT_RAM_3D = 256'h00F00FFFFFFFFFFFFFFFFFC000003FFFFFFFF00003FFFFFFFFFFFFFFFFF01F00;
defparam prom_inst_1.INIT_RAM_3E = 256'h00700FFFFFFFFFFFFFFFFFC000003FFFFFFFF00003FFFFFFFFFFFFFFFFF01E00;
defparam prom_inst_1.INIT_RAM_3F = 256'h00780FFFFFFFFFFFFFFFFFC000003FFFFFFFF00003FFFFFFFFFFFFFFFFF01E00;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h00780FFFFFFFFFFFFFFFFFF000003FFFFFFFF00003FFFFFFFFFFFFFFFFF01E00;
defparam prom_inst_2.INIT_RAM_01 = 256'h00780FFFFFFFFFFFFFFFFFF000003FFFFFFFF00003FFFFFFFFFFFFFFFFE01E00;
defparam prom_inst_2.INIT_RAM_02 = 256'h00780FFFFFFFFFFFFFFFFFF000003FFFFFFFF00003FFFFFFFFFFFFFFFFE01E00;
defparam prom_inst_2.INIT_RAM_03 = 256'h007807FFFFFFFFFFFFFFFFF000001FFFFFFFF00001FFFFFFFFFFFFFFFFE01E00;
defparam prom_inst_2.INIT_RAM_04 = 256'h007807FFFFFFFFFFFFFFFFF000001FFFFFFFF80001FFFFFFFFFFFFFFFFE01C00;
defparam prom_inst_2.INIT_RAM_05 = 256'h003C07FFFFFFFFFFFFFFFFF000001FFFFFFFF80001FFFFFFFFFFFFFFFFE03C00;
defparam prom_inst_2.INIT_RAM_06 = 256'h003C07FFFFFFFFFFFFFFFFF000001FFFFFFFF80001FFFFFFFFFFFFFFFFE03C00;
defparam prom_inst_2.INIT_RAM_07 = 256'h003C07FFFFFFFFFFFFFFFFF000001FFFFFFFF80000FFFFFFFFFFFFFFFFC03C00;
defparam prom_inst_2.INIT_RAM_08 = 256'h003C03FFFFFFFFFFFFFFFFF000001FFFFFFFF80000FFFFFFFFFFFFFFFFC03C00;
defparam prom_inst_2.INIT_RAM_09 = 256'h001C03FFFFFFFFFFFFFFFFF000001FFFFFFFF80000FFFFFFFFFFFFFFFFC03800;
defparam prom_inst_2.INIT_RAM_0A = 256'h001E03FFFFFFFFFFFFFFFFF000001FFFFFFFF800007FFFFFFFFFFFFFFFC07800;
defparam prom_inst_2.INIT_RAM_0B = 256'h001E03FFFFFFFFFFFFFFFFF000001FFFFFFFF800007FFFFFFFFFFFFFFFC07800;
defparam prom_inst_2.INIT_RAM_0C = 256'h001E01FFFFFFFFFFFFFFFFF000001FFFFFFFF800007FFFFFFFFFFFFFFF807800;
defparam prom_inst_2.INIT_RAM_0D = 256'h001E01FFFFFFFFFFFFFFFFF000001FFFFFFFF800003FFFFFFFFFFFFFFF807000;
defparam prom_inst_2.INIT_RAM_0E = 256'h000F81FFFFFFFFFFFFFFFFF000001FFFFFFFFC00003FFFFFFFFFFFFFFF81F000;
defparam prom_inst_2.INIT_RAM_0F = 256'h000F81FFFFFFFFFFFFFFFFF000001FFFFFFFFC00003FFFFFFFFFFFFFFF81F000;
defparam prom_inst_2.INIT_RAM_10 = 256'h000F81FFFFFFFFFFFFFFFFF000000FFFFFFFFC00003FFFFFFFFFFFFFFF81F000;
defparam prom_inst_2.INIT_RAM_11 = 256'h000F80FFFFFFFFFFFFFFFFF000000FFFFFFFFC00001FFFFFFFFFFFFFFF01F000;
defparam prom_inst_2.INIT_RAM_12 = 256'h000F80FFFFFFFFFFFFFFFFF000000FFFFFFFFC00001FFFFFFFFFFFFFFF01E000;
defparam prom_inst_2.INIT_RAM_13 = 256'h0007C0FFFFFFFFFFFFFFFFF000000FFFFFFFFC00001FFFFFFFFFFFFFFF03E000;
defparam prom_inst_2.INIT_RAM_14 = 256'h0007C0FFFFFFFFFFFFFFFFF000000FFFFFFFFC00000FFFFFFFFFFFFFFF03E000;
defparam prom_inst_2.INIT_RAM_15 = 256'h0007C07FFFFFFFFFFFFFFFF800000FFFFFFFFC00000FFFFFFFFFFFFFFE03E000;
defparam prom_inst_2.INIT_RAM_16 = 256'h0007C07FFFFFFFFFFFFFFFF800000FFFFFFFFC000007FFFFFFFFFFFFFE03C000;
defparam prom_inst_2.INIT_RAM_17 = 256'h0003E07FFFFFFFFFFFFFFFF800000FFFFFFFFC000007FFFFFFFFFFFFFE07C000;
defparam prom_inst_2.INIT_RAM_18 = 256'h0003C07FFFFFFFFFFFFFFFF800000FFFFFFFFE000007FFFFFFFFFFFFFE07C000;
defparam prom_inst_2.INIT_RAM_19 = 256'h0003E03FFFFFFFFFFFFFFFF800000FFFFFFFFE000003FFFFFFFFFFFFFC07C000;
defparam prom_inst_2.INIT_RAM_1A = 256'h0003E03FFFFFFFFFFFFFFFF800000FFFFFFFFE000003FFFFFFFFFFFFFC0F8000;
defparam prom_inst_2.INIT_RAM_1B = 256'h0003E03FFFFFFFFFFFFFFFF800000FFFFFFFFE000001FFFFFFFFFFFFFC0F8000;
defparam prom_inst_2.INIT_RAM_1C = 256'h0001F00FFFFFFFFFFFFFFFF8000007FFFFFFFE000001FFFFFFFFFFFFFC0F8000;
defparam prom_inst_2.INIT_RAM_1D = 256'h0001F00FFFFFFFFFFFFFFFF8000007FFFFFFFE000001FFFFFFFFFFFFFC0F8000;
defparam prom_inst_2.INIT_RAM_1E = 256'h0001F00FFFFFFFFFFFFFFFF0000007FFFFFFFE0000007FFFFFFFFFFFF00E0000;
defparam prom_inst_2.INIT_RAM_1F = 256'h0001F00FFFFFFFFFFFFFFFF0000007FFFFFFFE0000007FFFFFFFFFFFF01E0000;
defparam prom_inst_2.INIT_RAM_20 = 256'h0001F00FFFFFFFFFFFFFFFF0000007FFFFFFFF0000003FFFFFFFFFFFF01E0000;
defparam prom_inst_2.INIT_RAM_21 = 256'h00007807FFFFFFFFFFFFFFF0000007FFFFFFFF0000001FFFFFFFFFFFE01E0000;
defparam prom_inst_2.INIT_RAM_22 = 256'h00007807FFFFFFFFFFFFFFF0000007FFFFFFFF0000001FFFFFFFFFFFE01C0000;
defparam prom_inst_2.INIT_RAM_23 = 256'h00007807FFFFFFFFFFFFFFF0000007FFFFFFFF0000000FFFFFFFFFFFE03C0000;
defparam prom_inst_2.INIT_RAM_24 = 256'h00003C03FFFFFFFFFFFFFFF0000007FFFFFFFF0000000FFFFFFFFFFFE03C0000;
defparam prom_inst_2.INIT_RAM_25 = 256'h00003C03FFFFFFFFFFFFFFF0000007FFFFFFFF00000007FFFFFFFFFFC0380000;
defparam prom_inst_2.INIT_RAM_26 = 256'h00003C03FFFFC1FFFFFFFFF0000007FFFFFFFF00000007FFFFFFFFFFC0780000;
defparam prom_inst_2.INIT_RAM_27 = 256'h00001E01FFFFC1FFFFFFFFF0000007FFFFFFFF80000003FFFFFFFFFF80780000;
defparam prom_inst_2.INIT_RAM_28 = 256'h00001E01FFFFC1FFFFFFFFC0000007FFFFFFFF80000001FFFFFFFFFF80700000;
defparam prom_inst_2.INIT_RAM_29 = 256'h00001E01FFFFC0FFFFFFFFC0000007FFFFFFFF80000001FFFFFFFFFF80700000;
defparam prom_inst_2.INIT_RAM_2A = 256'h00001E01FFFFC0FFFFFFFFC0000007FFFFFFFF80000001FFFFFFFFFF80700000;
defparam prom_inst_2.INIT_RAM_2B = 256'h00000F00FFFFC0FFFFFFFFC0000007FFFFFFFF80000000FFFFFFFFFF00F00000;
defparam prom_inst_2.INIT_RAM_2C = 256'h00000F00FFFFE0FFFFFFFFC0000007FFFFFFFF800000007FFFFFFFFF00E00000;
defparam prom_inst_2.INIT_RAM_2D = 256'h00000F00FFFFE07FFFFFFFC0000007FFFFFFFFC00000007FFFFFFFFF00E00000;
defparam prom_inst_2.INIT_RAM_2E = 256'h000007807FFFE07FFFFFFF80000007FFFFFFFFC00000003FFFFFFFFE01E00000;
defparam prom_inst_2.INIT_RAM_2F = 256'h000007807FFFE07FFFFFFF80000007FFFFFFFFC00000000FFFFFFFFE01E00000;
defparam prom_inst_2.INIT_RAM_30 = 256'h000007807FFFE03FFFFFFF80000007FFFFFFFFC000000007FFFFFFFE03C00000;
defparam prom_inst_2.INIT_RAM_31 = 256'h000003C03FFFF00FFFFFFF00000007FFFFFFFFC000000007FFFFFFFC03C00000;
defparam prom_inst_2.INIT_RAM_32 = 256'h000003C03FFFF007FFFFFF00000007FFFFFFFFF000000003FFFFFFFC03C00000;
defparam prom_inst_2.INIT_RAM_33 = 256'h000003C03FFFF007FFFFFE00000007FFFFFFFFF000000001FFFFFFF80F800000;
defparam prom_inst_2.INIT_RAM_34 = 256'h000001F01FFFF803FFFFFE00000007FFFFFFFFF000000001FFFFFFF80F800000;
defparam prom_inst_2.INIT_RAM_35 = 256'h000001F01FFFF800FFFFFC00000007FFFFFFFFF000000000FFFFFFF80F800000;
defparam prom_inst_2.INIT_RAM_36 = 256'h000001F80FFFF8007FFFF800000007FFFFFFFFF800000000FFFFFFF01F000000;
defparam prom_inst_2.INIT_RAM_37 = 256'h000000F80FFFFC000FFFF000000007FFFFFFFFF8000000007FFFFFF01F000000;
defparam prom_inst_2.INIT_RAM_38 = 256'h000000F80FFFFC000FFFF000000007FFFFFFFFF8000000007FFFFFF01F000000;
defparam prom_inst_2.INIT_RAM_39 = 256'h000000F80FFFFC0001FF8000000007FFFFFFFFF8000000003FFFFFC01F000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h0000007C03FFFC0000000000000007FFFFFFFFF8000000003FFFFFC03E000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000007C03FFFE0000000000000007FFFFFFFFFC000000001FFFFFC03E000000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000007C01FFFE000000000000000FFFFFFFFFFC000000001FFFFF803C000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000003E01FFFF000000000000000FFFFFFFFFFC000000000FFFFF807C000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000003E00FFFF000000000000000FFFFFFFFFFC000000000FFFFF007C000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000000F00FFFF800000000000001FFFFFFFFFFE000000000FFFFF00F0000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0000000F007FFF800000000000001FFFFFFFFFFE000000000FFFFF00F0000000;
defparam prom_inst_3.INIT_RAM_01 = 256'h00000007807FFFC00000000000001FFFFFFFFFFE0000000003FFFE01E0000000;
defparam prom_inst_3.INIT_RAM_02 = 256'h00000007803FFFC00000000000003FFFFFFFFFFF0000000003FFFE01E0000000;
defparam prom_inst_3.INIT_RAM_03 = 256'h00000007803FFFF00000000000003FFFFFFFFFFF0000000003FFFC03C0000000;
defparam prom_inst_3.INIT_RAM_04 = 256'h00000003C03FFFF80000000000007FFFFFFFFFFF0000000003FFFC03C0000000;
defparam prom_inst_3.INIT_RAM_05 = 256'h00000003C01FFFF8000000000001FFFFFFFFFFFF800000000FFFF807C0000000;
defparam prom_inst_3.INIT_RAM_06 = 256'h00000003C01FFFF8000000000001FFFFFFFFFFFF800000000FFFF807C0000000;
defparam prom_inst_3.INIT_RAM_07 = 256'h00000001E01FFFFC000000000001FFFFFFFFFFFF800000000FFFF80780000000;
defparam prom_inst_3.INIT_RAM_08 = 256'h00000001E00FFFFE000000000003FFFFFFFFFFFFC00000000FFFF00780000000;
defparam prom_inst_3.INIT_RAM_09 = 256'h00000000F00FFFFF000000000007FFFFFFFFFFFFC00000000FFFF00F00000000;
defparam prom_inst_3.INIT_RAM_0A = 256'h00000000F007FFFF80000000000FFFFFFFFFFFFFE00000001FFFE00F00000000;
defparam prom_inst_3.INIT_RAM_0B = 256'h000000007C07FFFFC0000000001FFFFFFFFFFFFFF00000003FFFE03E00000000;
defparam prom_inst_3.INIT_RAM_0C = 256'h000000007C03FFFFF0000000003FFFFFFFFFFFFFFC0000003FFFC03E00000000;
defparam prom_inst_3.INIT_RAM_0D = 256'h000000003E03FFFFFC000000007FFFFFFFFFFFFFFE0000007FFFC07C00000000;
defparam prom_inst_3.INIT_RAM_0E = 256'h000000003E01FFFFFF00000000FFFFFFFFFFFFFFFF000000FFFF807C00000000;
defparam prom_inst_3.INIT_RAM_0F = 256'h000000001F007FFFFFC0000003FFFFFFFFFFFFFFFF800003FFFE00F800000000;
defparam prom_inst_3.INIT_RAM_10 = 256'h000000001F007FFFFFF000001FFFFFFFFFFFFFFFFFE00007FFFE01F800000000;
defparam prom_inst_3.INIT_RAM_11 = 256'h000000000F803FFFFFFF80007FFFFFFFFFFFFFFFFFF800FFFFFC01F000000000;
defparam prom_inst_3.INIT_RAM_12 = 256'h000000000F803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03F000000000;
defparam prom_inst_3.INIT_RAM_13 = 256'h000000000F803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03F000000000;
defparam prom_inst_3.INIT_RAM_14 = 256'h0000000003C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803C000000000;
defparam prom_inst_3.INIT_RAM_15 = 256'h0000000003E01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF807C000000000;
defparam prom_inst_3.INIT_RAM_16 = 256'h0000000001E00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0078000000000;
defparam prom_inst_3.INIT_RAM_17 = 256'h0000000001F007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00F8000000000;
defparam prom_inst_3.INIT_RAM_18 = 256'h0000000000F007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00F0000000000;
defparam prom_inst_3.INIT_RAM_19 = 256'h0000000000F803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01E0000000000;
defparam prom_inst_3.INIT_RAM_1A = 256'h00000000007801FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803E0000000000;
defparam prom_inst_3.INIT_RAM_1B = 256'h00000000003C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803C0000000000;
defparam prom_inst_3.INIT_RAM_1C = 256'h00000000003E00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00780000000000;
defparam prom_inst_3.INIT_RAM_1D = 256'h00000000001E007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00780000000000;
defparam prom_inst_3.INIT_RAM_1E = 256'h00000000001F807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01F00000000000;
defparam prom_inst_3.INIT_RAM_1F = 256'h00000000000FC03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03F00000000000;
defparam prom_inst_3.INIT_RAM_20 = 256'h000000000007C00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003E00000000000;
defparam prom_inst_3.INIT_RAM_21 = 256'h000000000007C00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003E00000000000;
defparam prom_inst_3.INIT_RAM_22 = 256'h000000000007E00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007C00000000000;
defparam prom_inst_3.INIT_RAM_23 = 256'h000000000003F007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00FC00000000000;
defparam prom_inst_3.INIT_RAM_24 = 256'h000000000001F003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01F800000000000;
defparam prom_inst_3.INIT_RAM_25 = 256'h000000000001F801FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF801E000000000000;
defparam prom_inst_3.INIT_RAM_26 = 256'h0000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF807E000000000000;
defparam prom_inst_3.INIT_RAM_27 = 256'h0000000000003C00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007C000000000000;
defparam prom_inst_3.INIT_RAM_28 = 256'h0000000000001E007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00F8000000000000;
defparam prom_inst_3.INIT_RAM_29 = 256'h0000000000001F003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00F8000000000000;
defparam prom_inst_3.INIT_RAM_2A = 256'h0000000000000F803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01F0000000000000;
defparam prom_inst_3.INIT_RAM_2B = 256'h00000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803E0000000000000;
defparam prom_inst_3.INIT_RAM_2C = 256'h00000000000007C00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003C0000000000000;
defparam prom_inst_3.INIT_RAM_2D = 256'h00000000000003F003FFFFFFFFFFFFFFFFFFFFFFFFFFFFC00F80000000000000;
defparam prom_inst_3.INIT_RAM_2E = 256'h00000000000001F801FFFFFFFFFFFFFFFFFFFFFFFFFFFF801F80000000000000;
defparam prom_inst_3.INIT_RAM_2F = 256'h00000000000001F801FFFFFFFFFFFFFFFFFFFFFFFFFFFF801F80000000000000;
defparam prom_inst_3.INIT_RAM_30 = 256'h00000000000000FC00FFFFFFFFFFFFFFFFFFFFFFFFFFFF003F00000000000000;
defparam prom_inst_3.INIT_RAM_31 = 256'h000000000000007E00FFFFFFFFFFFFFFFFFFFFFFFFFFFE007E00000000000000;
defparam prom_inst_3.INIT_RAM_32 = 256'h000000000000007E007FFFFFFFFFFFFFFFFFFFFFFFFFFE007C00000000000000;
defparam prom_inst_3.INIT_RAM_33 = 256'h000000000000003F003FFFFFFFFFFFFFFFFFFFFFFFFFFC00FC00000000000000;
defparam prom_inst_3.INIT_RAM_34 = 256'h000000000000000F801FFFFFFFFFFFFFFFFFFFFFFFFFF801F000000000000000;
defparam prom_inst_3.INIT_RAM_35 = 256'h0000000000000007C00FFFFFFFFFFFFFFFFFFFFFFFFFF003E000000000000000;
defparam prom_inst_3.INIT_RAM_36 = 256'h0000000000000003E007FFFFFFFFFFFFFFFFFFFFFFFFE007C000000000000000;
defparam prom_inst_3.INIT_RAM_37 = 256'h0000000000000003F003FFFFFFFFFFFFFFFFFFFFFFFFC00F8000000000000000;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000000000000001FC01FFFFFFFFFFFFFFFFFFFFFFFF803F0000000000000000;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000FC007FFFFFFFFFFFFFFFFFFFFFFE007E0000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h00000000000000007E003FFFFFFFFFFFFFFFFFFFFFFC00FE0000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h00000000000000003F001FFFFFFFFFFFFFFFFFFFFFF800FC0000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h00000000000000003F001FFFFFFFFFFFFFFFFFFFFFF800FC0000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h00000000000000001F800FFFFFFFFFFFFFFFFFFFFFF001F80000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h00000000000000000FC007FFFFFFFFFFFFFFFFFFFFE003F00000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h000000000000000003E003FFFFFFFFFFFFFFFFFFFF8007C00000000000000000;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h000000000000000003F001FFFFFFFFFFFFFFFFFFFF000F800000000000000000;
defparam prom_inst_4.INIT_RAM_01 = 256'h000000000000000001F8007FFFFFFFFFFFFFFFFFFE001F000000000000000000;
defparam prom_inst_4.INIT_RAM_02 = 256'h000000000000000000FC003FFFFFFFFFFFFFFFFFFC003E000000000000000000;
defparam prom_inst_4.INIT_RAM_03 = 256'h0000000000000000007E000FFFFFFFFFFFFFFFFFF0007C000000000000000000;
defparam prom_inst_4.INIT_RAM_04 = 256'h0000000000000000003F8007FFFFFFFFFFFFFFFFE001F8000000000000000000;
defparam prom_inst_4.INIT_RAM_05 = 256'h0000000000000000001FC003FFFFFFFFFFFFFFFF8007F0000000000000000000;
defparam prom_inst_4.INIT_RAM_06 = 256'h0000000000000000000FE000FFFFFFFFFFFFFFFF000FE0000000000000000000;
defparam prom_inst_4.INIT_RAM_07 = 256'h00000000000000000007F0007FFFFFFFFFFFFFFE001FC0000000000000000000;
defparam prom_inst_4.INIT_RAM_08 = 256'h00000000000000000001F8003FFFFFFFFFFFFFFC003F80000000000000000000;
defparam prom_inst_4.INIT_RAM_09 = 256'h000000000000000000007E000FFFFFFFFFFFFFF000FE00000000000000000000;
defparam prom_inst_4.INIT_RAM_0A = 256'h000000000000000000007E000FFFFFFFFFFFFFF000FE00000000000000000000;
defparam prom_inst_4.INIT_RAM_0B = 256'h000000000000000000003F0003FFFFFFFFFFFFC000FC00000000000000000000;
defparam prom_inst_4.INIT_RAM_0C = 256'h000000000000000000001F8001FFFFFFFFFFFF0001F800000000000000000000;
defparam prom_inst_4.INIT_RAM_0D = 256'h000000000000000000000FC0007FFFFFFFFFFE000FF000000000000000000000;
defparam prom_inst_4.INIT_RAM_0E = 256'h0000000000000000000007F0003FFFFFFFFFF8001FE000000000000000000000;
defparam prom_inst_4.INIT_RAM_0F = 256'h0000000000000000000003FC000FFFFFFFFFF0003FC000000000000000000000;
defparam prom_inst_4.INIT_RAM_10 = 256'h0000000000000000000001FE0007FFFFFFFFC0007F0000000000000000000000;
defparam prom_inst_4.INIT_RAM_11 = 256'h00000000000000000000007F0001FFFFFFFF8001FE0000000000000000000000;
defparam prom_inst_4.INIT_RAM_12 = 256'h00000000000000000000003FC0003FFFFFFC0003FC0000000000000000000000;
defparam prom_inst_4.INIT_RAM_13 = 256'h00000000000000000000000FE0001FFFFFF00007F00000000000000000000000;
defparam prom_inst_4.INIT_RAM_14 = 256'h000000000000000000000007F00007FFFFE0003FC00000000000000000000000;
defparam prom_inst_4.INIT_RAM_15 = 256'h000000000000000000000001FE0001FFFF80007F800000000000000000000000;
defparam prom_inst_4.INIT_RAM_16 = 256'h000000000000000000000000FF00007FFE0001FF000000000000000000000000;
defparam prom_inst_4.INIT_RAM_17 = 256'h0000000000000000000000007FC0003FF00003FC000000000000000000000000;
defparam prom_inst_4.INIT_RAM_18 = 256'h0000000000000000000000007FC0003FF00003FC000000000000000000000000;
defparam prom_inst_4.INIT_RAM_19 = 256'h0000000000000000000000001FE00007C0000FF8000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1A = 256'h0000000000000000000000000FF8000000001FF0000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1B = 256'h00000000000000000000000001FE000000007F80000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1C = 256'h00000000000000000000000000FF80000003FF00000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1D = 256'h000000000000000000000000003FE0000007FC00000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1E = 256'h000000000000000000000000001FF800001FF800000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1F = 256'h0000000000000000000000000007FE00007FE000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_20 = 256'h0000000000000000000000000001FF8001FF8000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_21 = 256'h00000000000000000000000000007FF00FFC0000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_22 = 256'h00000000000000000000000000001FFC3FF80000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_23 = 256'h000000000000000000000000000007FFFFE00000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_24 = 256'h000000000000000000000000000001FFFF800000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_25 = 256'h000000000000000000000000000001FFFF800000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_26 = 256'h0000000000000000000000000000007FFE000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_27 = 256'h0000000000000000000000000000000FF0000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_28 = 256'h00000000000000000000000000000003C0000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(dout[0]),
  .I0(mux_o_3),
  .I1(prom_inst_4_dout[0]),
  .S0(dff_q_0)
);
endmodule //logo_rom
