//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2AR-LV18EQ144C8/I7
//Device: GW2AR-18C
//Created Time: Mon Nov 07 09:50:32 2022

module cos_table (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h1F1E1D1C1B1A191817161514131211100F0E0D0C0B0A09080706050403020100;
defparam prom_inst_0.INIT_RAM_01 = 256'h3F3E3D3C3B3A393837363534333231302F2E2D2C2B2A29282726252423222120;
defparam prom_inst_0.INIT_RAM_02 = 256'h5F5E5D5C5B5A595857565554535251504F4E4D4C4B4A49484746454443424140;
defparam prom_inst_0.INIT_RAM_03 = 256'h7F7E7D7C7B7A797877767574737271706F6E6D6C6B6A69686766656463626160;
defparam prom_inst_0.INIT_RAM_04 = 256'h1F1E1D1C1A191817161514131211100F0E0D0C0B0A0908070605040302010000;
defparam prom_inst_0.INIT_RAM_05 = 256'h3F3E3D3C3B3A393837363534333231302F2E2D2C2B2A29282726252423222120;
defparam prom_inst_0.INIT_RAM_06 = 256'h5F5E5D5C5B5A595857565554535251504F4E4D4C4B4A49484746454443424140;
defparam prom_inst_0.INIT_RAM_07 = 256'h7F7E7D7C7B7A797877767574737271706F6E6D6C6B6A69686766656463626160;
defparam prom_inst_0.INIT_RAM_08 = 256'h1D1C1B1A191817161514131211100F0E0D0C0B0A090807060504030201000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h3E3D3C3B3A3938373635343332312F2E2D2C2B2A292827262524232221201F1E;
defparam prom_inst_0.INIT_RAM_0A = 256'h5E5D5C5B5A595857565554535251504F4E4D4C4B4A494847464544434241403F;
defparam prom_inst_0.INIT_RAM_0B = 256'h7F7E7D7C7B7A797877767574737271706F6E6D6C6B6A6968676664636261605F;
defparam prom_inst_0.INIT_RAM_0C = 256'h1B1A1918171514131211100F0E0D0C0B0A090807060504030201000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h3C3B3A393837363534333231302F2D2C2B2A292827262524232221201F1E1D1C;
defparam prom_inst_0.INIT_RAM_0E = 256'h5E5D5B5A595857565554535251504F4E4D4C4B4A4948474644434241403F3E3D;
defparam prom_inst_0.INIT_RAM_0F = 256'h7F7E7D7C7B7A7978777675747271706F6E6D6C6B6A696867666564636261605F;
defparam prom_inst_0.INIT_RAM_10 = 256'h17161514131211100E0D0C0B0A09080706050403010000000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h3A3938363534333231302F2E2D2C2B2A2827262524232221201F1E1D1B1A1918;
defparam prom_inst_0.INIT_RAM_12 = 256'h5C5B5A5958575655545352504F4E4D4C4B4A4948474645434241403F3E3D3C3B;
defparam prom_inst_0.INIT_RAM_13 = 256'h7F7E7D7C7B7A7977767574737271706F6E6D6C6A696867666564636261605F5D;
defparam prom_inst_0.INIT_RAM_14 = 256'h1211100F0E0C0B0A090807060503020100000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h363534333231302F2D2C2B2A2928272524232221201F1D1C1B1A191817161413;
defparam prom_inst_0.INIT_RAM_16 = 256'h5B5A58575655545352514F4E4D4C4B4A4947464544434241403E3D3C3B3A3938;
defparam prom_inst_0.INIT_RAM_17 = 256'h7F7E7D7C7A7978777675747371706F6E6D6C6B6968676665646362605F5E5D5C;
defparam prom_inst_0.INIT_RAM_18 = 256'h0B0A090807050403020100000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h3231302E2D2C2B2A28272625242221201F1E1C1B1A19181615141311100F0E0D;
defparam prom_inst_0.INIT_RAM_1A = 256'h58575655545251504F4E4C4B4A49484645444342403F3E3D3C3A393837363433;
defparam prom_inst_0.INIT_RAM_1B = 256'h7F7E7D7B7A79787775747372716F6E6D6C6B6968676665636261605F5D5C5B5A;
defparam prom_inst_0.INIT_RAM_1C = 256'h0302000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h2C2B2A282726242322211F1E1D1B1A19181615141211100E0D0C0B0908070504;
defparam prom_inst_0.INIT_RAM_1E = 256'h56545352504F4E4D4B4A49474645434241403E3D3C3A39383735343331302F2D;
defparam prom_inst_0.INIT_RAM_1F = 256'h7F7E7C7B7A797776757372716F6E6D6C6A69686665646361605F5D5C5B595857;
defparam prom_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h242322201F1D1C1B191816151412110F0E0C0B0A080705040301000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h52504F4D4C4B494846454442413F3E3D3B3A383735343331302E2D2C2A292726;
defparam prom_inst_0.INIT_RAM_23 = 256'h7F7E7C7B797877757472716F6E6D6B6A686766646361605E5D5C5A5957565553;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h1A1817151412110F0D0C0A090706040201000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_26 = 256'h4D4B494846454341403E3D3B3A3836353332302F2D2B2A2827252422201F1D1C;
defparam prom_inst_0.INIT_RAM_27 = 256'h7F7D7C7A7977767472716F6E6C6A6967666463615F5E5C5B595856545351504E;
defparam prom_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h0C0A080605030100000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2A = 256'h454442403E3C3B3937353332302E2C2A2927252321201E1C1A18171513110F0E;
defparam prom_inst_0.INIT_RAM_2B = 256'h7F7D7B7A78767472716F6D6B6968666462605F5D5B5957565452504E4D4B4947;
defparam prom_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2E = 256'h3B39373533302E2C2A282624221F1D1B19171513110E0C0A0806040200000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h7F7D7B79777472706E6C6A686663615F5D5B59575552504E4C4A484644413F3D;
defparam prom_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h2B292624211E1C191714110F0C0A070402000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h7F7C7A7775726F6D6A686562605D5A585553504D4B484643403E3B393633312E;
defparam prom_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h110D0A0603000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h7F7C7875716E6A6763605D5956524F4B4844413D3A3733302C2925221E1B1814;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h7F7A75706A65605B56514C47413C37322D28231E18130E090400000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h7F756B60564C42382D23190F0500000000000000000000000000000000000000;

endmodule //cos_table
