//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2AR-LV18EQ144C8/I7
//Device: GW2AR-18C
//Created Time: Fri Jun 02 19:02:27 2023

module table_FONT (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [16:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [0:0] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [0:0] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [0:0] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [0:0] prom_inst_7_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_0.INIT = 16'h0002;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_1.INIT = 16'h0008;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_2.INIT = 16'h0020;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_3.INIT = 16'h0080;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_4.INIT = 16'h0200;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_5.INIT = 16'h0800;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_6.INIT = 16'h2000;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_7.INIT = 16'h8000;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000020100000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000003E000001E0000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000010000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000C002000C0000000100000000000000000000000000000060000010;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000080040000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000010000000000008000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h000000000000000000000000000000000000000000001FC000F8000000000010;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000020100000000000000001000000000000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h0000000000000000002000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h0000000003E000001E000000000000000000000000000000000000007DE00000;
defparam prom_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000030000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000001C002000E0000000100000000000000000000000000000060000010;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000080040000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000000000000000000010000000000008000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000080040000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000010000000000008000000002000088000000000010;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h0010000000000000000000000060100000000000000002000000000000000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000000000000000006000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h00000000020020000200000000000000000000000000000000000000CFC00000;
defparam prom_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000020000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000000001000200020000000100000000000000000000000000000060000010;
defparam prom_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000080040000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h0000000000000000000000010000000000008000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000080040000000000000000;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000000000000000000000010000000000008000000002000188000000000010;
defparam prom_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h0010000000000000000000000040180000000000000002000440000000000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h0000000000000000006000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000F80;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000000002002000020000000000000000000000000000000000000000800000;
defparam prom_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000020000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000000003000200020000000200000000000000000000000000000060000010;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000080040000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000010000000000008000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000080040000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000010000000000008000000002000108000000000010;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h00200300000000000000000000C0080000000100000002000440000003000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h030000000000000000C0030000C0030000000400030000000300000000000300;
defparam prom_inst_1.INIT_RAM_04 = 256'h03000000000000000000018000000300060000000000000006000000000018C0;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000000002003000020000000000000000000000030000000300000003000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h0300000000000000000001800000000020000000070003000700060000000000;
defparam prom_inst_1.INIT_RAM_07 = 256'h0000000002000200020000000200000000000000018006000300000060000010;
defparam prom_inst_1.INIT_RAM_08 = 256'h0000030000000000000800000000000007000000000080040000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h0000180003800000000000010000000000008000000000000030000006000000;
defparam prom_inst_1.INIT_RAM_0A = 256'h00000300000000000018000000000000070000000700800400000000030000C0;
defparam prom_inst_1.INIT_RAM_0B = 256'h0000180003000000000000010000000000008000000006400108000007000010;
defparam prom_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_10 = 256'hF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FC0000;
defparam prom_inst_1.INIT_RAM_11 = 256'hF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FC;
defparam prom_inst_1.INIT_RAM_12 = 256'h00200780000000000000000000C00C00000037C01E000200044000000700F8FC;
defparam prom_inst_1.INIT_RAM_13 = 256'h078000000000000000C0078003E00FC001001F000FC03F000FC03FF83FF00F80;
defparam prom_inst_1.INIT_RAM_14 = 256'h0FC060FDF87EFFF9E0FC07E03FF00FC83FC007F87FFC0FF81F801FFDF87E1060;
defparam prom_inst_1.INIT_RAM_15 = 256'h000000000200100002003FF01FE0F87C303003000FC01FE00FC980FC0FC007F8;
defparam prom_inst_1.INIT_RAM_16 = 256'h0FC0F8FDC63EFFF9E0FC07E03FF0F8FC21803FF01FC1E7C01FC01F9DF87E0000;
defparam prom_inst_1.INIT_RAM_17 = 256'hF8FC00000200020002003FF00600F87C18600300E7C03F801FD01FF863000610;
defparam prom_inst_1.INIT_RAM_18 = 256'hF8FC0FC0F8FDF87EF83FE0F9F81DF81C1FE1878E7FFCFFFC07F81FFC1FFDF87E;
defparam prom_inst_1.INIT_RAM_19 = 256'hFC0E7E3E0FE01FFDF3FE3FE1FFFFFFFEFF00FFFCF87C0FC000781FE01F8007F8;
defparam prom_inst_1.INIT_RAM_1A = 256'hF8FC0FC0F8FDF87EF83CE0F8F81CF81C3FF1C78E1FC0FFFC07F81FF81FC0F3F0;
defparam prom_inst_1.INIT_RAM_1B = 256'h7C183E7E0FE00FF9F3FE3FC1FFFFFFFEFE00FFFCF87C3FE002001FE01FC00610;
defparam prom_inst_1.INIT_RAM_1C = 256'hF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FC;
defparam prom_inst_1.INIT_RAM_1D = 256'hF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FC;
defparam prom_inst_1.INIT_RAM_1E = 256'hF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FC;
defparam prom_inst_1.INIT_RAM_1F = 256'h0000F8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FCF8FC;
defparam prom_inst_1.INIT_RAM_20 = 256'hF878F878F878F878F878F878F878F878F878F878F878F878F878F878F8780000;
defparam prom_inst_1.INIT_RAM_21 = 256'hF878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878;
defparam prom_inst_1.INIT_RAM_22 = 256'h00200780000000000200000000800C000000346031000200044000000780F878;
defparam prom_inst_1.INIT_RAM_23 = 256'h078000080000400001C00780062018400300118018603E0018703FF83FF008C0;
defparam prom_inst_1.INIT_RAM_24 = 256'h18607079F03CFFF8E0F80C703FF0187860E007F87FF81FF830C03FF9F03C0020;
defparam prom_inst_1.INIT_RAM_25 = 256'h000000000200100002003FF01FE0F07C3030030018601FE01879C0F8186007F0;
defparam prom_inst_1.INIT_RAM_26 = 256'h18607079C61CFFF8E0F80C703FF0F87827E03FF07060EC60306030DDF03C0000;
defparam prom_inst_1.INIT_RAM_27 = 256'hF87800000200020002003FF00600F878186007006C6060C030701FF06FC01F90;
defparam prom_inst_1.INIT_RAM_28 = 256'h78781860F879F03CF826E0F8F83CF83C3039C78E7FF8FFFC03F83FF83FF9F03C;
defparam prom_inst_1.INIT_RAM_29 = 256'hFC0CC31C18303FF9F7FE7FE1FFFDFFFC7E00FFF8F07C078000881FE030C007F0;
defparam prom_inst_1.INIT_RAM_2A = 256'h787818607878F07CF864E0F8F83CF83C7038C78C7060FFFC03F83FF838607E10;
defparam prom_inst_1.INIT_RAM_2B = 256'h7C18633C18301FF1F7FCFFC1FFFCFFFC7E00FFFCF878233003001FE030601F90;
defparam prom_inst_1.INIT_RAM_2C = 256'hF878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878;
defparam prom_inst_1.INIT_RAM_2D = 256'hF878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878;
defparam prom_inst_1.INIT_RAM_2E = 256'hF878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878;
defparam prom_inst_1.INIT_RAM_30 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_1.INIT_RAM_31 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_1.INIT_RAM_32 = 256'h0040078000000000020000000180040000000C20210007900440000003002030;
defparam prom_inst_1.INIT_RAM_33 = 256'h078000180000600001C0078008001020020020C0103008001010201802001860;
defparam prom_inst_1.INIT_RAM_34 = 256'h3030701040088040203018100200203840300020403030206020601040080020;
defparam prom_inst_1.INIT_RAM_35 = 256'h0000000002001800020020100200601030700700102002002038403030300040;
defparam prom_inst_1.INIT_RAM_36 = 256'h303020304208804020301810020020302C200080403070306020207040080000;
defparam prom_inst_1.INIT_RAM_37 = 256'h20300000020002000200202005002030186005803820404020100080786030D0;
defparam prom_inst_1.INIT_RAM_38 = 256'h2010303020304008204620202030203060184208403020300040601060104008;
defparam prom_inst_1.INIT_RAM_39 = 256'h20088108101860104408C0404208420820002010601002000188020060200040;
defparam prom_inst_1.INIT_RAM_3A = 256'h20303030203043082044302020702070400842184030202000C0602020301808;
defparam prom_inst_1.INIT_RAM_3B = 256'h3030C118301830204408808042084208200010102030621807000200602030D0;
defparam prom_inst_1.INIT_RAM_3C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_1.INIT_RAM_3D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_1.INIT_RAM_3E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000203020302030203020302030203020302030203020302030203020302030;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_2.INIT_RAM_01 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_02 = 256'h004007800000000002000000018004000000082020801FD00440000000002030;
defparam prom_inst_2.INIT_RAM_03 = 256'h000000700000300001C007801800303002002040301008002000003002001020;
defparam prom_inst_2.INIT_RAM_04 = 256'h201070104008804020301008020020184010002040306020C030401040080010;
defparam prom_inst_2.INIT_RAM_05 = 256'h0000000002000800020020300200203030500580203002002018603020100040;
defparam prom_inst_2.INIT_RAM_06 = 256'h2010203042088040203010080200203038100080001070104010603040080000;
defparam prom_inst_2.INIT_RAM_07 = 256'h2030000002000200020020600D00102018E00480303000402010008070302070;
defparam prom_inst_2.INIT_RAM_08 = 256'h2010201020304008204630202070207040044208403020200040401040104008;
defparam prom_inst_2.INIT_RAM_09 = 256'h201081882008401048088040420842082000201020300F8001080200C0300040;
defparam prom_inst_2.INIT_RAM_0A = 256'h20302010203043082044102020502050400022100010204000C0402060101008;
defparam prom_inst_2.INIT_RAM_0B = 256'h3020811820082020440880804208420820001010102042080500020040102070;
defparam prom_inst_2.INIT_RAM_0C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_0D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_0E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_0F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_10 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_2.INIT_RAM_11 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_12 = 256'h0040000000000000020000000180060000001C30208010300440000000002030;
defparam prom_inst_2.INIT_RAM_13 = 256'h000000C000001C00038000003000201002006040200008002000006002003020;
defparam prom_inst_2.INIT_RAM_14 = 256'h6018681040088040303010080200601840180020403040204010C01060100010;
defparam prom_inst_2.INIT_RAM_15 = 256'h0000000002000800020020200200102028500480201002006018203060180040;
defparam prom_inst_2.INIT_RAM_16 = 256'h4018203042088040303010080200203030180080001860080010403060100000;
defparam prom_inst_2.INIT_RAM_17 = 256'h2030000002000200020020C0090018602CA00480203000402010008070184030;
defparam prom_inst_2.INIT_RAM_18 = 256'h2010601820304008204210202050205040006210403020600040C010C0106010;
defparam prom_inst_2.INIT_RAM_19 = 256'h201180882008C01048098040420842082000201010201FE00108020040100040;
defparam prom_inst_2.INIT_RAM_1A = 256'h20304018203045082040182020D020D0400022100018204000C0402040181008;
defparam prom_inst_2.INIT_RAM_1B = 256'h30608098600020204C0880804208420820001010186042080580020000104030;
defparam prom_inst_2.INIT_RAM_1C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_1D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_1E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_1F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_20 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_2.INIT_RAM_21 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_22 = 256'h00800000000000000200000001000600000014102080303004C0000000002030;
defparam prom_inst_2.INIT_RAM_23 = 256'h0000018000000600038000002000201006004020200008002000004002002030;
defparam prom_inst_2.INIT_RAM_24 = 256'h4008681040088040103010080200401840080020403040200018801020100010;
defparam prom_inst_2.INIT_RAM_25 = 256'h0000000002000C00020020600200186028500480201002004018303040080040;
defparam prom_inst_2.INIT_RAM_26 = 256'h4008203042088040103010080200203030080080000860080018401020100000;
defparam prom_inst_2.INIT_RAM_27 = 256'h20300000020002000200008008800CC024B008C0203000402000008060084010;
defparam prom_inst_2.INIT_RAM_28 = 256'h2010400820304008204010202050205040002210403020400040801080102010;
defparam prom_inst_2.INIT_RAM_29 = 256'h2031008840008010480900404208420820002010186032300300020000180040;
defparam prom_inst_2.INIT_RAM_2A = 256'h20304008203044882040082020902090400032200008204000C0402040081008;
defparam prom_inst_2.INIT_RAM_2B = 256'h30C1809840002020440880804208420821C010100CC042080C80020000184010;
defparam prom_inst_2.INIT_RAM_2C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_2D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_2E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_2F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_30 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_2.INIT_RAM_31 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_32 = 256'h00800000000000000200000001000600000016302100201004C0000000002030;
defparam prom_inst_2.INIT_RAM_33 = 256'h0000030000000300000000002000201004004020200008006000008002002010;
defparam prom_inst_2.INIT_RAM_34 = 256'h40086C1040088040103010080200400040080020403080200008801020103E10;
defparam prom_inst_2.INIT_RAM_35 = 256'h0000000002000400020020400200084028500880201002004000103040080040;
defparam prom_inst_2.INIT_RAM_36 = 256'h4008203042088040103010080200203020080080000860080008C01020100000;
defparam prom_inst_2.INIT_RAM_37 = 256'h2030000002000200020001801880048024900840203000402000008060084010;
defparam prom_inst_2.INIT_RAM_38 = 256'h2010400820304008204018202090209040002210403020400040801080102010;
defparam prom_inst_2.INIT_RAM_39 = 256'h2021008840008010480900404208420820002010084062180300020000080040;
defparam prom_inst_2.INIT_RAM_3A = 256'h20304008203044882040042021902190600012200008204000C06020C0081018;
defparam prom_inst_2.INIT_RAM_3B = 256'h3F8100984000202044088080420842082FE010100480C20808C0020000084010;
defparam prom_inst_2.INIT_RAM_3C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_3D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_3E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000203020302030203020302030203020302030203020302030203020302030;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_3.INIT_RAM_01 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_02 = 256'h0080000000000000020000000100060000001220110020103FF8000000002030;
defparam prom_inst_3.INIT_RAM_03 = 256'h02000E00FFF8018000000000200020100400402060003FF02000018002002010;
defparam prom_inst_3.INIT_RAM_04 = 256'hC008641043088040183010080200600040080020003080200008C0103FF01310;
defparam prom_inst_3.INIT_RAM_05 = 256'h0000000002000400020020C002000CC068D008402010020060001830C0080040;
defparam prom_inst_3.INIT_RAM_06 = 256'h400820304208804018301008020020302008008000086008000880103FF00000;
defparam prom_inst_3.INIT_RAM_07 = 256'h203000000200020001000100108007002590084020300040180000806008C010;
defparam prom_inst_3.INIT_RAM_08 = 256'h2010C00820304308204008202090209040002230003020400040C010C0103FF0;
defparam prom_inst_3.INIT_RAM_09 = 256'h206100884000C010480980404208420821C020100CC042080300020000080040;
defparam prom_inst_3.INIT_RAM_0A = 256'h2030400820304C8820400620211021103E001A400008204040C03020C0081030;
defparam prom_inst_3.INIT_RAM_0B = 256'h3FC100987F8018204708E080420842083C3010100700C208084002000008C010;
defparam prom_inst_3.INIT_RAM_0C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_0D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_0E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_0F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_10 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_3.INIT_RAM_11 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_12 = 256'h01000000000000000200000001000600000033201E0820003FF0000002002030;
defparam prom_inst_3.INIT_RAM_13 = 256'h02001800FFFC00E0000000004000203004004060200008102000030002002010;
defparam prom_inst_3.INIT_RAM_14 = 256'h800C6410430880400830100802002000FE080C2006308020000840103FE01110;
defparam prom_inst_3.INIT_RAM_15 = 256'h000000000200060002000080020004804C9008402010020020000C30800C0040;
defparam prom_inst_3.INIT_RAM_16 = 256'h40082030420880400830100802002030200800807FF86008000880103FE00000;
defparam prom_inst_3.INIT_RAM_17 = 256'h20301C000E000200018002001040030027101040203000400F80008060088010;
defparam prom_inst_3.INIT_RAM_18 = 256'h2010800C2030430820400C202190219060001220063020400040401040103FE0;
defparam prom_inst_3.INIT_RAM_19 = 256'h20C10088C00040104C0880404208420827E020100480C2080500020000080040;
defparam prom_inst_3.INIT_RAM_1A = 256'h203040083FF04848204003E0221022100FC00FC07FF8204040C01FE0C0081FE0;
defparam prom_inst_3.INIT_RAM_1B = 256'h306100F87F800FE043F87F8042084208301010100300C2081040420800088010;
defparam prom_inst_3.INIT_RAM_1C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_1D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_1E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_1F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_20 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_3.INIT_RAM_21 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_22 = 256'h0100000000000000020000000100060000002160003020000480000002002030;
defparam prom_inst_3.INIT_RAM_23 = 256'h0200300000000030000000004780302004006060200008302000020002002010;
defparam prom_inst_3.INIT_RAM_24 = 256'h800C6210450800400C30100802003000FC080C20063080200008601010201110;
defparam prom_inst_3.INIT_RAM_25 = 256'h00000000020002000200018002000700449818402010020030000630800C1FC0;
defparam prom_inst_3.INIT_RAM_26 = 256'h40082030420800400C3010080200203020080080400860080008C01010200000;
defparam prom_inst_3.INIT_RAM_27 = 256'h20303E080C00020001C0060030400700231010202030004001E000806008C010;
defparam prom_inst_3.INIT_RAM_28 = 256'h2010800C20304508204004202110211030001260063020400040601060101020;
defparam prom_inst_3.INIT_RAM_29 = 256'h21810088C00060104408C040420842082C3020100700820C0580020000081FC0;
defparam prom_inst_3.INIT_RAM_2A = 256'h2030400820304848204003202610261038000EC04008204040C01FE0C0081FC0;
defparam prom_inst_3.INIT_RAM_2B = 256'h30210098400000204008008042084208201010100700C208106042080008C010;
defparam prom_inst_3.INIT_RAM_2C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_2D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_2E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_2F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_3.INIT_RAM_30 = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF00000;
defparam prom_inst_3.INIT_RAM_31 = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_3.INIT_RAM_32 = 256'h010000007FF800007FF8084001000600000001C000E030000480000003003FF0;
defparam prom_inst_3.INIT_RAM_33 = 256'h0600E0000000001C000000004DC018600C0020E0200008201000060002002010;
defparam prom_inst_3.INIT_RAM_34 = 256'h80046210458800400670100002001E0000080FE007F0802000083FF010201110;
defparam prom_inst_3.INIT_RAM_35 = 256'h0000000002000200020001000300030044981060201002001E0007F080043840;
defparam prom_inst_3.INIT_RAM_36 = 256'h40082030420800400670100002003FF020080080400860084018401010200000;
defparam prom_inst_3.INIT_RAM_37 = 256'h3FF0221002000200010004002060048063101020203000400020008060084010;
defparam prom_inst_3.INIT_RAM_38 = 256'h201080043FF0458820400620231023101FC01A4007F0204000403FF03FF01020;
defparam prom_inst_3.INIT_RAM_39 = 256'h3F8100F8FF803FF047F87FC04208420838102010030082040C80020000083840;
defparam prom_inst_3.INIT_RAM_3A = 256'h2030400820305848204006202410241060080A404008204040C0302040081000;
defparam prom_inst_3.INIT_RAM_3B = 256'h3021809840080020400800844208420820101010048042083020420840184010;
defparam prom_inst_3.INIT_RAM_3C = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_3.INIT_RAM_3D = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_3.INIT_RAM_3E = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_3.INIT_RAM_3F = 256'h00003FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF00000;
defparam prom_inst_4.INIT_RAM_01 = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_4.INIT_RAM_02 = 256'h020000007FF800007FF808C0010006000000008003001C000480000003003FF0;
defparam prom_inst_4.INIT_RAM_03 = 256'h0C006000000000180300030058400FC0080030A02000082018000C0002002010;
defparam prom_inst_4.INIT_RAM_04 = 256'h800463104488004003F01000020007C000080FE007F0802000080FF010601110;
defparam prom_inst_4.INIT_RAM_05 = 256'h00000000020003000200030003000300448810202010020007C01C3080046040;
defparam prom_inst_4.INIT_RAM_06 = 256'h401820304208004003F0100002003FF030080080600860084010403010600000;
defparam prom_inst_4.INIT_RAM_07 = 256'h3FF061300200020003000C10202008C043183020203000402030018060084010;
defparam prom_inst_4.INIT_RAM_08 = 256'h201080043FF04488204003E0221022100FC00FC007F0204000400FF01FF01060;
defparam prom_inst_4.INIT_RAM_09 = 256'h20E100F8FF801FF041F83FC04208420830102010030082040880020000086040;
defparam prom_inst_4.INIT_RAM_0A = 256'h2030401820305028204044202C102C10401012206008204040C0202040181000;
defparam prom_inst_4.INIT_RAM_0B = 256'h302080982008002040080084420842082010101008C042082020420840104010;
defparam prom_inst_4.INIT_RAM_0C = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_4.INIT_RAM_0D = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_4.INIT_RAM_0E = 256'h3FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_4.INIT_RAM_0F = 256'h00003FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF03FF0;
defparam prom_inst_4.INIT_RAM_10 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_4.INIT_RAM_11 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_12 = 256'h02000000000002000200048001000600020000800C0007800480000003002030;
defparam prom_inst_4.INIT_RAM_13 = 256'h10003800000000700780078050600FC008001FA0302008400F00080002002010;
defparam prom_inst_4.INIT_RAM_14 = 256'h800C61104C88004001B010000200006000080C20063080200008181008401110;
defparam prom_inst_4.INIT_RAM_15 = 256'h00000000020001000200020005800700448810202010020000603030800C4040;
defparam prom_inst_4.INIT_RAM_16 = 256'h201020304208004001B010000200203030180080201870106010603008400000;
defparam prom_inst_4.INIT_RAM_17 = 256'h203001E002000200020018304020186040082010203000402010038070184030;
defparam prom_inst_4.INIT_RAM_18 = 256'h2010800C20304C88204003A02210221018000EC0063020400040181000100840;
defparam prom_inst_4.INIT_RAM_19 = 256'h20210088C00000104008004042084208201020100700820C08C0020000084040;
defparam prom_inst_4.INIT_RAM_1A = 256'h203020102030502820404C2028102810401092242018204040C0202060181000;
defparam prom_inst_4.INIT_RAM_1B = 256'h3020811820180020400800844208420820101010186042082010420860104030;
defparam prom_inst_4.INIT_RAM_1C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_1D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_1E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_1F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_20 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_4.INIT_RAM_21 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_22 = 256'h02000000000003000200058001800600030000C0300000C00C80000003002030;
defparam prom_inst_4.INIT_RAM_23 = 256'h30000C00FFFC00C0078007806020186008000E2018E008400F00100002002010;
defparam prom_inst_4.INIT_RAM_24 = 256'h8008619048C80040013010000200002000080C20063080200008201008401310;
defparam prom_inst_4.INIT_RAM_25 = 256'h0000000002000100020006000480048047083020201002000020203080084040;
defparam prom_inst_4.INIT_RAM_26 = 256'h3030307047180040013010000200203038100080303070306020207008400000;
defparam prom_inst_4.INIT_RAM_27 = 256'h2030004002000200020010304030302040082010203000403030868070102070;
defparam prom_inst_4.INIT_RAM_28 = 256'h20108008203048C8204002202410241020000A40063020408040201000100840;
defparam prom_inst_4.INIT_RAM_29 = 256'h20110088400000104008004242084208201020100480C2081040020000084040;
defparam prom_inst_4.INIT_RAM_2A = 256'h203030302030702820404820381038106030A2343030204040C0302020381000;
defparam prom_inst_4.INIT_RAM_2B = 256'h3020C11830180020400800844208420820101010302062184010420860202070;
defparam prom_inst_4.INIT_RAM_2C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_2D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_2E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_2F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_30 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_4.INIT_RAM_31 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_32 = 256'h040000000000030002000300018004000300004041C000207FF0218003002030;
defparam prom_inst_4.INIT_RAM_33 = 256'h20000600000001800780078060201020180000200FA008C01800100002002010;
defparam prom_inst_4.INIT_RAM_34 = 256'hC008609048480040023010000200001000080420023080200008201008401E10;
defparam prom_inst_4.INIT_RAM_35 = 256'h00002010020001800200040008C00C80430820302010420800102030C0088040;
defparam prom_inst_4.INIT_RAM_36 = 256'h186018F8453C00400230100002002030EC303FE018606C60706030D008400000;
defparam prom_inst_4.INIT_RAM_37 = 256'h203000000200020002003FF1E0707878F03CF87C38381FF83860CCF0F86030DC;
defparam prom_inst_4.INIT_RAM_38 = 256'h2010C00820304848204006202410241060081A40023020408040201000100840;
defparam prom_inst_4.INIT_RAM_39 = 256'h20110088400000104008004242084208201020100C8042081060420800088040;
defparam prom_inst_4.INIT_RAM_3A = 256'h7FF818607078E01C7FE070F8F07CF07C3070E71C18607FE07FF01FF838681870;
defparam prom_inst_4.INIT_RAM_3B = 256'h7FE0633818780071F01C03FCE33CE33C7878383878782330E03C7FF8706030DC;
defparam prom_inst_4.INIT_RAM_3C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_3D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_3E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_4.INIT_RAM_3F = 256'h0000203020302030203020302030203020302030203020302030203020302030;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_5.INIT_RAM_01 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_02 = 256'h0400000000000300020003000180040003000040022000200880308003002030;
defparam prom_inst_5.INIT_RAM_03 = 256'h2000030000000700030003006020302010000020002008803000200002002010;
defparam prom_inst_5.INIT_RAM_04 = 256'h40086090584800400630100002000010000880202030C0204008201008C01C10;
defparam prom_inst_5.INIT_RAM_05 = 256'h0000303002000080020008100840084043082010201042080010603040088040;
defparam prom_inst_5.INIT_RAM_06 = 256'h0FC00FB83DEE00400630100002002030E7E03FF00FC067C05FC01F9008C00000;
defparam prom_inst_5.INIT_RAM_07 = 256'h203000000200020002003FF0F0787878F03CF87C3C3C3FF82FC078F1EFC01F9C;
defparam prom_inst_5.INIT_RAM_08 = 256'h2010400820305848204004202C102C10400812202030204080402010201008C0;
defparam prom_inst_5.INIT_RAM_09 = 256'h2011008840080010400800424208420820102010084062183020420840088040;
defparam prom_inst_5.INIT_RAM_0A = 256'h7FF80FC07879E01CFFF070F8E07CE07C1FD0C78C0FC0FFF07FF80FF81FC80FE0;
defparam prom_inst_5.INIT_RAM_0B = 256'h7FC03E7C0FE800F9F03E03FDE79DE79CFC7C787C78783FE1F07C7FF85FC01F9C;
defparam prom_inst_5.INIT_RAM_0C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_0D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_0E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_0F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_10 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_5.INIT_RAM_11 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_12 = 256'h040000000000030002000FC000800C000300004002100020088030C003002030;
defparam prom_inst_5.INIT_RAM_13 = 256'h200001C000000C00000000002020203010000020002008802000200002002010;
defparam prom_inst_5.INIT_RAM_14 = 256'h40186050506800400C3010000200201040188020603040204018601004801010;
defparam prom_inst_5.INIT_RAM_15 = 256'h000010200200008002000810106018604308201020104208201020304018C040;
defparam prom_inst_5.INIT_RAM_16 = 256'h0300060010C000400C3010000200203001800080030063000700061004800000;
defparam prom_inst_5.INIT_RAM_17 = 256'h2030000002000200020000000000000000000000000000400300000003000600;
defparam prom_inst_5.INIT_RAM_18 = 256'h201040182030506820400C202810281040181220603020408040601060100480;
defparam prom_inst_5.INIT_RAM_19 = 256'h201100884008001040080042420842082010201018603A70202042084018C040;
defparam prom_inst_5.INIT_RAM_1A = 256'h0000030000000000000000000000000007080000030000000000000003080300;
defparam prom_inst_5.INIT_RAM_1B = 256'h000018000300000000000000000000000000000000000A400000000007000600;
defparam prom_inst_5.INIT_RAM_1C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_1D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_1E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_1F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_20 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_5.INIT_RAM_21 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_22 = 256'h080000000000030002003B7000800C00030004C004101020088030C003002030;
defparam prom_inst_5.INIT_RAM_23 = 256'h2020006000001800000000002020201010000040002009002000201002002030;
defparam prom_inst_5.INIT_RAM_24 = 256'h6010605050280040183010000200201040108020603040204010201004801010;
defparam prom_inst_5.INIT_RAM_25 = 256'h00001840020000C0020010101020102040084010201042082010203060104040;
defparam prom_inst_5.INIT_RAM_26 = 256'h0000000000000040183010000200203000000080000060000000001004800000;
defparam prom_inst_5.INIT_RAM_27 = 256'h2030000002000200020000000000000000000000000000400000000000000000;
defparam prom_inst_5.INIT_RAM_28 = 256'h2010601020305028204088203810381040193234603020408040201060100480;
defparam prom_inst_5.INIT_RAM_29 = 256'h201180886008001040080042420842082010201010201FE02030420840104040;
defparam prom_inst_5.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000180000;
defparam prom_inst_5.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000002000000000000000000;
defparam prom_inst_5.INIT_RAM_2C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_2D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_2E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_2F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_30 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_5.INIT_RAM_31 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_32 = 256'h08000000000003000200231000C0080003000F8004103020088018E003002030;
defparam prom_inst_5.INIT_RAM_33 = 256'h3020003000003000000000002020203010000040002009002000201002003020;
defparam prom_inst_5.INIT_RAM_34 = 256'h2030607070280040103010000200203040308020603020206030201004801030;
defparam prom_inst_5.INIT_RAM_35 = 256'h000008C002000040020010103030303040084008201042082030303020304040;
defparam prom_inst_5.INIT_RAM_36 = 256'h0000000000000040103010000200203000000080000060000000001004800000;
defparam prom_inst_5.INIT_RAM_37 = 256'h2030000002000200020000000000000000000000000000400000000000000000;
defparam prom_inst_5.INIT_RAM_38 = 256'h2010203020307028204098203010301060192214603020408040201060100480;
defparam prom_inst_5.INIT_RAM_39 = 256'h2030810820180010400800424208420820102010303002006010420860304040;
defparam prom_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000780000000000000000000000000000000300000;
defparam prom_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000002000000000000000000;
defparam prom_inst_5.INIT_RAM_3C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_3D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_3E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_5.INIT_RAM_3F = 256'h0000203020302030203020302030203020302030203020302030203020302030;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h2030203020302030203020302030203020302030203020302030203020300000;
defparam prom_inst_6.INIT_RAM_01 = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_6.INIT_RAM_02 = 256'h0800000000000300020003000040080003000F00041030600880186003002030;
defparam prom_inst_6.INIT_RAM_03 = 256'h102000180000600000000000302030203010008000200B002000301002001020;
defparam prom_inst_6.INIT_RAM_04 = 256'h3020603060280040203010000200302060608020603030207020301007001020;
defparam prom_inst_6.INIT_RAM_05 = 256'h0000048002000040020020102010201040084008201042083020103030202040;
defparam prom_inst_6.INIT_RAM_06 = 256'h0000000000000040203010000200203000000180000060000000001007000400;
defparam prom_inst_6.INIT_RAM_07 = 256'h2030000002000200020000000000000000000000000000400000000000000000;
defparam prom_inst_6.INIT_RAM_08 = 256'h2010302020306028204090203010301030396214603020408040301060100700;
defparam prom_inst_6.INIT_RAM_09 = 256'h2060C30830380010400800424208420820102010201002004018420870202040;
defparam prom_inst_6.INIT_RAM_0A = 256'h0000000000000000000000000DC000000000000000000000000000000FE00000;
defparam prom_inst_6.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000002000000000000000000;
defparam prom_inst_6.INIT_RAM_0C = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_6.INIT_RAM_0D = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_6.INIT_RAM_0E = 256'h2030203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_6.INIT_RAM_0F = 256'h0000203020302030203020302030203020302030203020302030203020302030;
defparam prom_inst_6.INIT_RAM_10 = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F80000;
defparam prom_inst_6.INIT_RAM_11 = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_12 = 256'h100000000000070000000300004018000700000004103CC008801C60030078F8;
defparam prom_inst_6.INIT_RAM_13 = 256'h1CE000000000000000000000106010202010018000200A001030103002301060;
defparam prom_inst_6.INIT_RAM_14 = 256'h1CC0F83DE01C07F8F8FDFF803FF03CE078C0FFF87FFC1FF85CC01FFC03F01020;
defparam prom_inst_6.INIT_RAM_15 = 256'h000005800200006002003FF0F87CF87DF87FF87EF8FC7FF83CE01FFC1CC03FF8;
defparam prom_inst_6.INIT_RAM_16 = 256'h00000000000007F8F8FDFF803FF078F800000100000060000000001003F00600;
defparam prom_inst_6.INIT_RAM_17 = 256'h78F8000003000200020000000000000000000000000000400000000000000000;
defparam prom_inst_6.INIT_RAM_18 = 256'hFFFC1CC078F9E01CFFF0F0F9E0FDE0FC18C9C78C7FFCFFF0FFF81FFC7FFC03F0;
defparam prom_inst_6.INIT_RAM_19 = 256'hFFC0663E1CE800FDF07E03FFF7BFF7BEFC7CFCFCF87C0FC1F07C7FF85CC03FF8;
defparam prom_inst_6.INIT_RAM_1A = 256'h000000000000000000000000186000000000000000000000000000001FC00000;
defparam prom_inst_6.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000002000000000000000000;
defparam prom_inst_6.INIT_RAM_1C = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_1D = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_1E = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_1F = 256'h000078F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_20 = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F80000;
defparam prom_inst_6.INIT_RAM_21 = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_22 = 256'h100000000000070000000300006010000700000002201F8008800C70030078F8;
defparam prom_inst_6.INIT_RAM_23 = 256'h0FC00000000000000000000018C018602010030000200A001860186003E01840;
defparam prom_inst_6.INIT_RAM_24 = 256'h0780F81DE01C03F8F8FDFF803FF02F804F80FFF87FFC07F84F8007FC03F01840;
defparam prom_inst_6.INIT_RAM_25 = 256'h000003000200002002003FF0F07CF07CF87DF07EF87C7FF82F8007FC07800FF0;
defparam prom_inst_6.INIT_RAM_26 = 256'h00000000000003F8F8FDFF803FF078F80000C300000060000000001003F00300;
defparam prom_inst_6.INIT_RAM_27 = 256'h78F8000001000200060000000000000000000000000000400000000000000000;
defparam prom_inst_6.INIT_RAM_28 = 256'hFFFC078078F9E01CFFF0E0F8E07CE07C0F8887847FFCFFF0FFF807FC7FFC03F0;
defparam prom_inst_6.INIT_RAM_29 = 256'hFF803C3E0FC800FDF03E01FEE7BEE7BEF87CF87CF07C0781F03C7FF84F800FF0;
defparam prom_inst_6.INIT_RAM_2A = 256'h0000000000000000000000001020000000000000000000000000000030000000;
defparam prom_inst_6.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000003C00000000000000000;
defparam prom_inst_6.INIT_RAM_2C = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_2D = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_2E = 256'h78F878F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_2F = 256'h000078F878F878F878F878F878F878F878F878F878F878F878F878F878F878F8;
defparam prom_inst_6.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_32 = 256'h10000000000007800000030000201000078000000360020008800E3803000000;
defparam prom_inst_6.INIT_RAM_33 = 256'h0000000000000000000000000F800FC03FF07E001FE00C000FC00FC003800FC0;
defparam prom_inst_6.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000FC0;
defparam prom_inst_6.INIT_RAM_35 = 256'h0000030003E000201E0000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_36 = 256'h000000000000000000000000000000000000FE00000078000000001C00000100;
defparam prom_inst_6.INIT_RAM_37 = 256'h0000000001C002000C0000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3A = 256'h0000000000000000000000001020000000000000000000000000000020000000;
defparam prom_inst_6.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000003C00000000000000000;
defparam prom_inst_6.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_02 = 256'h2000000000000000000000000000000000000000008002000880000003000000;
defparam prom_inst_7.INIT_RAM_03 = 256'h0000000000000000000000000700070000003800000000000780078002000700;
defparam prom_inst_7.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000780;
defparam prom_inst_7.INIT_RAM_05 = 256'h0000010000000030000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000180;
defparam prom_inst_7.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_12 = 256'h2000000000000000000000000000000000000000000002000880000000000000;
defparam prom_inst_7.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_15 = 256'h0000000000000010000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000080;
defparam prom_inst_7.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_18 = 256'h0000000000000000000000000780000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_22 = 256'h2000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_25 = 256'h0000000000000010000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_28 = 256'h0000000000000000000000000DC0000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_38 = 256'h0000000000000000000000001860000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(prom_inst_4_dout[0]),
  .I1(prom_inst_5_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(prom_inst_6_dout[0]),
  .I1(prom_inst_7_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_1)
);
MUX2 mux_inst_6 (
  .O(dout[0]),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_0)
);
endmodule //table_FONT
