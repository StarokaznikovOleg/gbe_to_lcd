//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-3
//Part Number: GW2AR-LV18EQ144C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Fri Oct 06 21:03:57 2023

module bme240_i2cmem (dout, clk, oce, ce, reset, ad);

output [8:0] dout;
input clk;
input oce;
input ce;
input reset;
input [8:0] ad;

wire [26:0] promx9_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROMX9 promx9_inst_0 (
    .DO({promx9_inst_0_dout_w[26:0],dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,gw_gnd,ad[8:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_0.READ_MODE = 1'b0;
defparam promx9_inst_0.BIT_WIDTH = 9;
defparam promx9_inst_0.RESET_MODE = "SYNC";
defparam promx9_inst_0.INIT_RAM_00 = 288'h287D3E40013BD1DDF1FF863E9F200BC9DDF1FFFFFFFFFFFFFC21F4F97C1DFF1F9341DDF1;
defparam promx9_inst_0.INIT_RAM_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_02 = 288'hFFFFFFFFFFFFFD01F4F97C1DFF1F93CDDDF1000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_04 = 288'hF97C1DFF1F93E9DDF1F97C1DFF1F93E5DDF1F97C1DFF1F93E1DDF1F97C1DFF1F93DDDDF1;
defparam promx9_inst_0.INIT_RAM_05 = 288'hF97C1DFF1F93F9DDF1F97C1DFF1F93F5DDF1F97C1DFF1F93F1DDF1F97C1DFF1F93EDDDF1;
defparam promx9_inst_0.INIT_RAM_06 = 288'h0000000000000000000000000000000000000000000000000000000000000000000001F4;
defparam promx9_inst_0.INIT_RAM_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;
defparam promx9_inst_0.INIT_RAM_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000;

endmodule //bme240_i2cmem
