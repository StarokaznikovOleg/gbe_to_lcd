//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2AR-LV18EQ144C8/I7
//Device: GW2AR-18C
//Created Time: Tue Aug 29 17:49:31 2023

module table_TEXT (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h8C0092858288908F000000000000A5A8ADA5B9A1AEAEB100A5AEB2B1A592232B;
defparam prom_inst_0.INIT_RAM_01 = 256'h25262400000000000000000000303000A0AAAEB0B29100003030000000219088;
defparam prom_inst_0.INIT_RAM_02 = 256'h8C0092858288908F000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h00262400000000000000000000313000A0AAAEB0B29100003130000000219088;
defparam prom_inst_0.INIT_RAM_04 = 256'h8C0092858288908F000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h00262400000000000000000000323000A0AAAEB0B29100003230000000219088;
defparam prom_inst_0.INIT_RAM_06 = 256'h8C0092858288908F000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h00262400000000000000000000333000A0AAAEB0B29100003330000000219088;
defparam prom_inst_0.INIT_RAM_08 = 256'h8C0092858288908F000000000000A5A8ADA5B9A1AEAEB100A5AEB2B1A592232A;
defparam prom_inst_0.INIT_RAM_09 = 256'h26252400000000000000000000303000A0AAAEB0B29100003430000000219088;
defparam prom_inst_0.INIT_RAM_0A = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_0B = 256'hF600000000000000000000000000000000000000000000003530000000219088;
defparam prom_inst_0.INIT_RAM_0C = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_0D = 256'hF600000000000000000000000000000000000000000000003630000000219088;
defparam prom_inst_0.INIT_RAM_0E = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_0F = 256'hF600000000000000000000000000000000000000000000003730000000219088;
defparam prom_inst_0.INIT_RAM_10 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_11 = 256'hF600000000000000000000000000000000000000000000003830000000219088;
defparam prom_inst_0.INIT_RAM_12 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_13 = 256'hF600000000000000000000000000000000000000000000003930000000219088;
defparam prom_inst_0.INIT_RAM_14 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_15 = 256'hF600000000000000000000000000000000000000000000003031000000219088;
defparam prom_inst_0.INIT_RAM_16 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_17 = 256'hF600000000000000000000000000000000000000000000003131000000219088;
defparam prom_inst_0.INIT_RAM_18 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_19 = 256'hF600000000000000000000000000000000000000000000003231000000219088;
defparam prom_inst_0.INIT_RAM_1A = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_1B = 256'hF600000000000000000000000000000000000000000000003331000000219088;
defparam prom_inst_0.INIT_RAM_1C = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_1D = 256'hF600000000000000000000000000000000000000000000003431000000219088;
defparam prom_inst_0.INIT_RAM_1E = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_1F = 256'hF600000000000000000000000000000000000000000000003531000000219088;
defparam prom_inst_0.INIT_RAM_20 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_21 = 256'hF600000000000000000000000000000000000000000000003631000000219088;
defparam prom_inst_0.INIT_RAM_22 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_23 = 256'hF600000000000000000000000000000000000000000000003731000000219088;
defparam prom_inst_0.INIT_RAM_24 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_25 = 256'hF600000000000000000000000000000000000000000000003831000000219088;
defparam prom_inst_0.INIT_RAM_26 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_27 = 256'hF600000000000000000000000000000000000000000000003931000000219088;
defparam prom_inst_0.INIT_RAM_28 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_29 = 256'hF600000000000000000000000000000000000000000000003032000000219088;
defparam prom_inst_0.INIT_RAM_2A = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_2B = 256'hF600000000000000000000000000000000000000000000003132000000219088;
defparam prom_inst_0.INIT_RAM_2C = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_2D = 256'hF600000000000000000000000000000000000000000000003232000000219088;
defparam prom_inst_0.INIT_RAM_2E = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_2F = 256'hF600000000000000000000000000000000000000000000003332000000219088;
defparam prom_inst_0.INIT_RAM_30 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_31 = 256'hF600000000000000000000000000000000000000000000003432000000219088;
defparam prom_inst_0.INIT_RAM_32 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_33 = 256'hF600000000000000000000000000000000000000000000003532000000219088;
defparam prom_inst_0.INIT_RAM_34 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_35 = 256'hF600000000000000000000000000000000000000000000003632000000219088;
defparam prom_inst_0.INIT_RAM_36 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_37 = 256'hF600000000000000000000000000000000000000000000003732000000219088;
defparam prom_inst_0.INIT_RAM_38 = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_39 = 256'hF600000000000000000000000000000000000000000000003832000000219088;
defparam prom_inst_0.INIT_RAM_3A = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_3B = 256'hF600000000000000000000000000000000000000000000003932000000219088;
defparam prom_inst_0.INIT_RAM_3C = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_3D = 256'hF600000000000000000000000000000000000000000000003033000000219088;
defparam prom_inst_0.INIT_RAM_3E = 256'h8C0092858288908F0000000000000000000000000000000000000000000000F6;
defparam prom_inst_0.INIT_RAM_3F = 256'hF600000000000000000000000000000000000000000000003133000000219088;

endmodule //table_TEXT
