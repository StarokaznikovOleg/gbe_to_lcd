//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-3
//Part Number: GW2AR-LV18EQ144C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Mon Nov 13 16:58:30 2023

module indexDDR_table (dout, clk, oce, ce, reset, ad);

output [11:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [19:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[19:0],dout[11:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h005A0054004E00480042003C00360030002A0024001E00180012000C00060000;
defparam prom_inst_0.INIT_RAM_01 = 256'h00BA00B400AE00A800A2009C00960090008A0084007E00780072006C00660060;
defparam prom_inst_0.INIT_RAM_02 = 256'h011A0114010E0108010200FC00F600F000EA00E400DE00D800D200CC00C600C0;
defparam prom_inst_0.INIT_RAM_03 = 256'h017A0174016E01680162015C01560150014A0144013E01380132012C01260120;
defparam prom_inst_0.INIT_RAM_04 = 256'h01DA01D401CE01C801C201BC01B601B001AA01A4019E01980192018C01860180;
defparam prom_inst_0.INIT_RAM_05 = 256'h023A0234022E02280222021C02160210020A020401FE01F801F201EC01E601E0;
defparam prom_inst_0.INIT_RAM_06 = 256'h029A0294028E02880282027C02760270026A0264025E02580252024C02460240;
defparam prom_inst_0.INIT_RAM_07 = 256'h02FA02F402EE02E802E202DC02D602D002CA02C402BE02B802B202AC02A602A0;
defparam prom_inst_0.INIT_RAM_08 = 256'h035A0354034E03480342033C03360330032A0324031E03180312030C03060300;
defparam prom_inst_0.INIT_RAM_09 = 256'h03BA03B403AE03A803A2039C03960390038A0384037E03780372036C03660360;
defparam prom_inst_0.INIT_RAM_0A = 256'h041A0414040E0408040203FC03F603F003EA03E403DE03D803D203CC03C603C0;
defparam prom_inst_0.INIT_RAM_0B = 256'h047A0474046E04680462045C04560450044A0444043E04380432042C04260420;
defparam prom_inst_0.INIT_RAM_0C = 256'h04DA04D404CE04C804C204BC04B604B004AA04A4049E04980492048C04860480;
defparam prom_inst_0.INIT_RAM_0D = 256'h053A0534052E05280522051C05160510050A050404FE04F804F204EC04E604E0;
defparam prom_inst_0.INIT_RAM_0E = 256'h059A0594058E05880582057C05760570056A0564055E05580552054C05460540;
defparam prom_inst_0.INIT_RAM_0F = 256'h05FA05F405EE05E805E205DC05D605D005CA05C405BE05B805B205AC05A605A0;
defparam prom_inst_0.INIT_RAM_10 = 256'h065A0654064E06480642063C06360630062A0624061E06180612060C06060600;
defparam prom_inst_0.INIT_RAM_11 = 256'h06BA06B406AE06A806A2069C06960690068A0684067E06780672066C06660660;
defparam prom_inst_0.INIT_RAM_12 = 256'h071A0714070E0708070206FC06F606F006EA06E406DE06D806D206CC06C606C0;
defparam prom_inst_0.INIT_RAM_13 = 256'h077A0774076E07680762075C07560750074A0744073E07380732072C07260720;
defparam prom_inst_0.INIT_RAM_14 = 256'h07DA07D407CE07C807C207BC07B607B007AA07A4079E07980792078C07860780;
defparam prom_inst_0.INIT_RAM_15 = 256'h083A0834082E08280822081C08160810080A080407FE07F807F207EC07E607E0;
defparam prom_inst_0.INIT_RAM_16 = 256'h089A0894088E08880882087C08760870086A0864085E08580852084C08460840;
defparam prom_inst_0.INIT_RAM_17 = 256'h08FA08F408EE08E808E208DC08D608D008CA08C408BE08B808B208AC08A608A0;
defparam prom_inst_0.INIT_RAM_18 = 256'h095A0954094E09480942093C09360930092A0924091E09180912090C09060900;
defparam prom_inst_0.INIT_RAM_19 = 256'h09BA09B409AE09A809A2099C09960990098A0984097E09780972096C09660960;
defparam prom_inst_0.INIT_RAM_1A = 256'h0A1A0A140A0E0A080A0209FC09F609F009EA09E409DE09D809D209CC09C609C0;
defparam prom_inst_0.INIT_RAM_1B = 256'h0A7A0A740A6E0A680A620A5C0A560A500A4A0A440A3E0A380A320A2C0A260A20;
defparam prom_inst_0.INIT_RAM_1C = 256'h0ADA0AD40ACE0AC80AC20ABC0AB60AB00AAA0AA40A9E0A980A920A8C0A860A80;
defparam prom_inst_0.INIT_RAM_1D = 256'h0B3A0B340B2E0B280B220B1C0B160B100B0A0B040AFE0AF80AF20AEC0AE60AE0;
defparam prom_inst_0.INIT_RAM_1E = 256'h0B9A0B940B8E0B880B820B7C0B760B700B6A0B640B5E0B580B520B4C0B460B40;
defparam prom_inst_0.INIT_RAM_1F = 256'h0BFA0BF40BEE0BE80BE20BDC0BD60BD00BCA0BC40BBE0BB80BB20BAC0BA60BA0;
defparam prom_inst_0.INIT_RAM_20 = 256'h0C5A0C540C4E0C480C420C3C0C360C300C2A0C240C1E0C180C120C0C0C060C00;
defparam prom_inst_0.INIT_RAM_21 = 256'h0CBA0CB40CAE0CA80CA20C9C0C960C900C8A0C840C7E0C780C720C6C0C660C60;
defparam prom_inst_0.INIT_RAM_22 = 256'h0D1A0D140D0E0D080D020CFC0CF60CF00CEA0CE40CDE0CD80CD20CCC0CC60CC0;
defparam prom_inst_0.INIT_RAM_23 = 256'h0D7A0D740D6E0D680D620D5C0D560D500D4A0D440D3E0D380D320D2C0D260D20;
defparam prom_inst_0.INIT_RAM_24 = 256'h0DDA0DD40DCE0DC80DC20DBC0DB60DB00DAA0DA40D9E0D980D920D8C0D860D80;
defparam prom_inst_0.INIT_RAM_25 = 256'h0E3A0E340E2E0E280E220E1C0E160E100E0A0E040DFE0DF80DF20DEC0DE60DE0;
defparam prom_inst_0.INIT_RAM_26 = 256'h0E9A0E940E8E0E880E820E7C0E760E700E6A0E640E5E0E580E520E4C0E460E40;
defparam prom_inst_0.INIT_RAM_27 = 256'h0EFA0EF40EEE0EE80EE20EDC0ED60ED00ECA0EC40EBE0EB80EB20EAC0EA60EA0;
defparam prom_inst_0.INIT_RAM_28 = 256'h0F5A0F540F4E0F480F420F3C0F360F300F2A0F240F1E0F180F120F0C0F060F00;
defparam prom_inst_0.INIT_RAM_29 = 256'h0FBA0FB40FAE0FA80FA20F9C0F960F900F8A0F840F7E0F780F720F6C0F660F60;
defparam prom_inst_0.INIT_RAM_2A = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FEA0FE40FDE0FD80FD20FCC0FC60FC0;
defparam prom_inst_0.INIT_RAM_2B = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_2C = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_2D = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_2E = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_2F = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_30 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_31 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_32 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_33 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_34 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_35 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_36 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_37 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_38 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_39 = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_3A = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_3B = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_3C = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_3D = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_3E = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;
defparam prom_inst_0.INIT_RAM_3F = 256'h0FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0;

endmodule //indexDDR_table
